
module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] anyedge
);
reg [7:0] prev_in;

always @(posedge clk) begin
  prev_in <= in;
  anyedge <= in ^ prev_in;   // 1 when any bit changes
end

endmodule
