
module TopModule (
    input clk,
    input load,
    input [511:0] data,
    output reg [511:0] q
);

  // Internal wire to hold the next state of the system
  wire [511:0] next_q;

  always @(posedge clk) begin
    if (load) begin
      // Load the current state with input data
      q <= data;
    end else begin
      // Advance by one time step using Rule 90 logic for each cell
      q[0] <= 0; // Left boundary is always 0
      q[511] <= 0; // Right boundary is always 0

      integer i;
      for (i = 1; i < 511; i = i + 1) begin
        next_q[i] = q[i-1] ^ q[i+1]; // Calculate the next state using Rule 90
      end

      // Update the current state with the next state
      for (i = 0; i <= 511; i = i + 1) begin
        if (!load) begin
          q[i] <= next_q[i];
        end
      end
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
