
module TopModule (
    input  wire [3:0] in,
    output wire [2:0] out_both,
    output wire [3:1] out_any,
    output wire [3:0] out_different
);

    /* 1) out_both[i] = in[i] & in[i+1]   (i = 2,1,0) */
    assign out_both[2] = in[2] & in[3];
    assign out_both[1] = in[1] & in[2];
    assign out_both[0] = in[0

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
