
module TopModule (
  output zero
);
  
  // Assign 0 to the output 'zero'
  zero = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
