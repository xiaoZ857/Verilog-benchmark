
module TopModule (
  input clk,
  input reset,
  input in,
  output reg disc,
  output reg flag,
  output reg err
);

  // State encoding
  typedef enum logic [2:0] {
    S0 = 3'b000, // Initial/default state
    S1 = 3'b001, // One consecutive '1'
    S2 = 3'b010, // Two consecutive '1's
    S3 = 3'b011, // Three consecutive '1's
    S4 = 3'b100, // Four consecutive '1's
    S5 = 3'b101, // Five consecutive '1's
    S6 = 3'b110, // Six consecutive '1's
    S7 = 3'b111  // Error state for seven or more consecutive '1's
  } state_t;

  state_t current_state, next_state;

  always_ff @(posedge clk or posedge reset) begin
    if (reset)
      current_state <= S0;
    else
      current_state <= next_state;
  end

  always_comb begin
    // Default output signals
    disc = 1'b0;
    flag = 1'b0;
    err = 1'b0;

    case (current_state)
      S0: begin
        if (in == 1'b1) 
          next_state = S1; 
        else 
          next_state = S0;
      end

      S1: begin
        if (in == 1'b1) 
          next_state = S2; 
        else 
          next_state = S0;
      end
      
      S2: begin
        if (in == 1'b1) 
          next_state = S3; 
        else 
          next_state = S0;
      end

      S3: begin
        if (in == 1'b1) 
          next_state = S4; 
        else 
          next_state = S0;
      end

      S4: begin
        if (in == 1'b1) 
          next_state = S5; 
        else 
          next_state = S0;
      end

      S5: begin
        if (in == 1'b1) 
          next_state = S6; 
        else begin
          // Discard the bit as it is a stuffed zero
          disc = 1'b1;
          next_state = S0;
        end
      end

      S6: begin
        if (in == 1'b1) 
          next_state = S7; 
        else begin
          // Detected flag sequence
          flag = 1'b1;
          next_state = S0;
        end
      end
      
      S7: begin
        err = 1'b1;
        next_state = S7; // Remain in error state for seven or more consecutive '1's
      end

    endcase
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
