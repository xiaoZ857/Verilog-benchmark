
module TopModule (
  input [3:0] in,
  output reg [1:0] pos
);
always @* begin
  if (in[0])          pos = 2'b00; // bit 0 is the first set bit
  else if (in[1])     pos = 2'b01; // bit 1 is the first set bit
  else if (in[2])     pos = 2'b10; // bit 2 is the first set bit
  else if (in[3])     pos = 2'b11; // bit 3 is the first set bit
  else                pos = 2'b00; // no bits set → output zero
end

endmodule
