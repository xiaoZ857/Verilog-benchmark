

module TopModule (
  input ring,
  input vibrate_mode,
  output ringer,
  output motor
);

always @(posedge clk) begin
    if (ring) begin
        if (vibrate_mode) begin
            ringer <= 0;
            motor <= 1;
        end else begin
            ringer <= 1;
            motor <= 0;
        end
    end else begin
        ringer <= 0;
        motor <= 0;
    end
end

endmodule
