
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
always @(posedge clk or posedge reset) begin
    if(reset) begin
        state <= 4'b0001; // Resetting to initial state A
    end else begin
        case (state)
            4'b0001: begin // State A
                if (w) state <= 4'b0010; // Transition to B on w=1
                else state <= 4'b0001; // Stay in A if w=0
            end,
            4'b0010: begin // State B
                if (!w) state <= 4'b0001; // Transition to A on w=0
                else if (w) state <= 4'b0011; // Stay in B or transition to D on w=1
            end,
            4'b0011: begin // State D
                if (!w) state <= 4'b1110; // Transition to A on w=0
                else if (w) state <= 4'b0111; // Stay in D or transition to E/C on w=1
            end,
            4'b0111: begin // State E (or C)
                if (!w) state <= 4'b0110; // Transition to D on w=0
                else state <= 4'b0111; // Stay in E or transition to D on w=1
            end,
            4'b1110: begin // State F
                if (w) state <= 4'b0100; // Transition to C on w=1
                else state <= 4'b1110; // Stay in F or transition to D on w=0
            end,
            4'b1111: begin // State A again (or D)
                if (w) state <= 4'b0010; // Transition to B on w=1
                else state <= 4'b1111; // Stay in A or transition to D on w=0
            enddefault: state <= 4'b0001; // Default state is A
        endcase
    end
end

always_comb begin
    z = (state == 4'b1110);
end

// VERILOG-EVAL: endmodule not found
