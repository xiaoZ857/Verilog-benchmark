
module TopModule (
    input clk,
    input j,
    input k,
    input areset,
    output reg out
);

    // State encoding
    typedef enum logic [1:0] {
        OFF = 2'b00,
        ON  = 2'b01
    } state_t;

    state_t current_state, next_state;

    // Output logic based on the current state
    always @(*) begin
        case (current_state)
            OFF: out = 1'b0;
            ON : out = 1'b1;
            default: out = 1'b0; // Default assignment to avoid latches
        endcase
    end

    // Next state logic and state register update
    always @(posedge clk or posedge areset) begin
        if (areset) begin
            current_state <= OFF;
        end else begin
            current_state <= next_state;
        end
    end

    // Next state logic based on the current state and inputs
    always @(*) begin
        case (current_state)
            OFF: 
                if (j == 1'b1) 
                    next_state = ON;  
                else 
                    next_state = OFF;

            ON: 
                if (k == 1'b1) 
                    next_state = OFF;
                else 
                    next_state = ON;

            default: 
                next_state = OFF;
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
