
module TopModule (
  input mode,
  input too_cold,
  input too_hot,
  input fan_on,
  output heater,
  output aircon,
  output fan
);
  // Heater is on only in heating mode when too_cold is asserted
  assign heater = mode & too_cold;
  
  // Air conditioner is on only in cooling mode when too_hot is asserted
  assign aircon = ~mode & too_hot;
  
  // Fan is on when either heater, air conditioner, or user request is active
  assign fan = heater | aircon | fan_on;

endmodule
