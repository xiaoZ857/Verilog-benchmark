
module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] pedge
);
reg [7:0] pedge_0;
reg [7:0] pedge_1;
reg [7:0] pedge_2;
reg [7:0] pedge_3;
reg [7:0] pedge_4;
reg [7:0] pedge_5;
reg [7:0] pedge_6;
reg [7:0] pedge_7;

always @(posedge clk) begin
  // Update the output bits based on the current input values
  if (in[0] == 0 && in[1] == 1) pedge_0 <= 1;
  else if (in[0] == 1 && in[1] == 0) pedge_0 <= 0;

  if (in[1] == 0 && in[2] == 1) pedge_1 <= 1;
  else if (in[1] == 1 && in[2] == 0) pedge_1 <= 0;

  if (in[2] == 0 && in[3] == 1) pedge_2 <= 1;
  else if (in[2] == 1 && in[3] == 0) pedge_2 <= 0;

  if (in[3] == 0 && in[4] == 1) pedge_3 <= 1;
  else if (in[3] == 1 && in[4] == 0) pedge_3 <= 0;

  if (in[4] == 0 && in[5] == 1) pedge_4 <= 1;
  else if (in[4] == 1 && in[5] == 0) pedge_4 <= 0;

  if (in[5] == 0 && in[6] == 1) pedge_5 <= 1;
  else if (in[5] == 1 && in[6] == 0) pedge_5 <= 0;

  if (in[6] == 0 && in[7] == 1) pedge_6 <= 1;
  else if (in[6] == 1 && in[7] == 0) pedge_6 <= 0;

  if (in[7] == 0 && in[0] == 1) pedge_7 <= 1;
  else if (in[7] == 1 && in[0] == 0) pedge_7 <= 0;

  // Assign the output bits to the main output
  pedge = {pedge_0, pedge_1, pedge_2, pedge_3, pedge_4, pedge_5, pedge_6, pedge_7};
end

endmodule
