
module TopModule (
  input clk,
  input shift_ena,
  input count_ena,
  input data,
  output reg [3:0] q
);

  always @(posedge clk) begin
    if (shift_ena) begin
      // Shift operation: insert new data at MSB, right-shift other bits
      q <= {data, q[3:1]};
    end else if (count_ena) begin
      // Down counter operation: decrement the current value
      q <= q - 4'b0001;
      
      // Handle wrap-around if the result is negative
      if (q == 4'b1111) begin
        q <= 4'b1110; // Wrap around to 14 when going below 0
      end
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
