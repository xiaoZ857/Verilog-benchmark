

module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);



// VERILOG-EVAL: endmodule not found
