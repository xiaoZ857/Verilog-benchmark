
module TopModule (
    input in,
    input [3:0] state,
    output reg [3:0] next_state,
    output out
);

// Output logic
assign out = (state == 4'b1000) ? 1 : 0;

always @(*) begin
    // Default to zero when no condition matches
    next_state = 4'b0000;

    case (state)
        4'b0001: // State A
            next_state = (!in) ? 4'b0001 : 4'b0010;
        4'b0010: // State B
            next_state = (!in) ? 4'b0100 : 4'b0010;
        4'b0100: // State C
            next_state = (!in) ? 4'b0001 : 4'b1000;
        4'b1000: // State D
            next_state = (!in) ? 4'b0100 : 4'b0010;
    endcase
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
