
module TopModule (
  input [4:1] x,
  output logic f
);
assign f = (~x[1] & ~x[2] & ~x[3] & ~x[4]) |  // 0000
           (~x[1] & ~x[2] & x[3] & ~x[4]) |   // 0010  
           (x[1] & x[2] & ~x[3] & ~x[4]) |    // 1100
           (x[1] & x[2] & ~x[3] & x[4]) |     // 1101
           (x[1] & x[2] & x[3] & x[4]) |      // 1111
           (x[1] & ~x[2] & ~x[3] & ~x[4]) |   // 1000
           (x[1] & ~x[2] & ~x[3] & x[4]) |    // 1001
           (x[1] & ~x[2] & x[3] & ~x[4]);     // 1010

endmodule
