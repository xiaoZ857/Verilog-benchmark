
module TopModule (
  input clk,
  input in,
  input reset,
  output done
);
  reg [2:0] state, next_state;
  reg [3:0] bit_count, next_bit_count;
  
  localparam IDLE = 3'b000;
  localparam START = 3'b001;
  localparam DATA  = 3'b010;
  localparam STOP  = 3'b011;
  localparam ERROR = 3'b100;
  
  always @(posedge clk) begin
    if (reset) begin
      state <= IDLE;
      bit_count <= 0;
    end else begin
      state <= next_state;
      bit_count <= next_bit_count;
    end
  end
  
  always @(*) begin
    next_state = state;
    next_bit_count = bit_count;
    
    case (state)
      IDLE: begin
        next_bit_count = 0;
        if (in == 1'b0) begin
          next_state = START;
        end
      end
      
      START: begin
        next_state = DATA;
        next_bit_count = 0;
      end
      
      DATA: begin
        if (bit_count == 7) begin
          next_state = STOP;
          next_bit_count = 0;
        end else begin
          next_bit_count = bit_count + 1;
        end
      end
      
      STOP: begin
        if (in == 1'b1) begin
          next_state = IDLE;
        end else begin
          next_state = ERROR;
        end
      end
      
      ERROR: begin
        if (in == 1'b1) begin
          next_state = IDLE;
        end
      end
      
      default: begin
        next_state = IDLE;
      end
    endcase
  end
  
  assign done = (state == STOP && in == 1'b1);
endmodule
