
module TopModule (
  input clk,
  input resetn,
  input x,
  input y,
  output f,
  output g
);
  // State definition
  typedef enum logic [1:0] {
    STATE_A,
    STATE_F_SET,
    STATE_X_MONITOR,
    STATE_G_SET,
    STATE_Y_MONITOR_1,
    STATE_Y_MONITOR_2
  } state_t;

  state_t current_state, next_state;

  // Registers for x history
  logic [2:0] x_history;

  // Registers for y monitoring
  logic [1:0] y_monitor_count;

  // Output registers
  logic f_reg, g_reg;

  // Assign outputs
  assign f = f_reg;
  assign g = g_reg;

  // State register update
  always_ff @(posedge clk, negedge resetn) begin
    if (!resetn) begin
      current_state <= STATE_A;
    end else begin
      current_state <= next_state;
    end
  end

  // Output register update
  always_ff @(posedge clk, negedge resetn) begin
    if (!resetn) begin
      f_reg <= 0;
      g_reg <= 0;
    end else begin
      case (current_state)
        STATE_F_SET: f_reg <= 1;
        STATE_G_SET: g_reg <= 1;
        default: ;
      endcase
    end
  end

  // Next state logic
  always_comb begin
    next_state = current_state;

    case (current_state)
      STATE_A: begin
        if (!resetn) begin
          next_state = STATE_A;
        end else begin
          next_state = STATE_F_SET;
        end
      end

      STATE_F_SET: begin
        next_state = STATE_X_MONITOR;
      end

      STATE_X_MONITOR: begin
        if (x) begin
          x_history[0] = 1;
        end else begin
          x_history[0] = 0;
        end

        if (x_history[0] == 1 && x_history[1] == 0 && x_history[2] == 1) begin
          next_state = STATE_G_SET;
        end else begin
          next_state = STATE_X_MONITOR;
        end
      end

      STATE_G_SET: begin
        y_monitor_count[0] = 0;
        y_monitor_count[1] = 0;
        next_state = STATE_Y_MONITOR_1;
      end

      STATE_Y_MONITOR_1: begin
        if (y) begin
          next_state = STATE_Y_MONITOR_2;
        end else begin
          y_monitor_count[0] = y_monitor_count[1];
          y_monitor_count[1] = 0;
          next_state = STATE_Y_MONITOR_1;
        end
      end

      STATE_Y_MONITOR_2: begin
        if (y) begin
          next_state = STATE_X_MONITOR;
        end else begin
          if (y_monitor_count[0] == 0 && y_monitor_count[1] == 0) begin
            next_state = STATE_Y_MONITOR_2;
          end else begin
            next_state = STATE_X_MONITOR;
          end
        end
      end

      default: begin
        next_state = STATE_A;
      end
    endcase
  end

  // Shift x history
  always_ff @(posedge clk, negedge resetn) begin
    if (!resetn) begin
      x_history[1:0] <= 0;
      x_history[2] <= 0;
    end else begin
      x_history[1:0] <= x_history[0:1];
      x_history[2] <= x_history[0];
    end
  end

endmodule
