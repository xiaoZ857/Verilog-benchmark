
module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);
reg [1:0] state, next_state;
assign out = (state == 2'b10);

always @(posedge clk or posedge reset) begin
    if (reset)
        state <= 2'b00;
    else
        state <= next_state;
end

always @(*) begin
    case(state)
        2'b00: if (j) next_state = 2'b10; else next_state = 2'b00;
        2'b10: if (~k) next_state = 2'b10; else next_state = 2'b00;
        default: next_state = 2'b00;
    endcase
end

endmodule
