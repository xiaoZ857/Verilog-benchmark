
module TopModule (
  input [7:0] in,
  output [31:0] out
);


// VERILOG-EVAL: endmodule not found
