
module TopModule (
  input in1,
  input in2,
  output logic out
);

// Implementing a 2-input NOR gate using the negation of OR operation
assign out = !(in1 | in2);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
