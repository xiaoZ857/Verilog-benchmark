
module TopModule (
  input clk,
  input d,
  output reg q
);
reg q;

always @(posedge clk) begin // Clocked by the positive edge of the clock signal
  if (d == 1) begin // If the data is high, set the output to 1
    q <= 1;
  else if (d == 0) begin // If the data is low, set the output to 0
    q <= 0;
  end
end

initial begin
  q = 0; // Default value of the flip-flop
end

// VERILOG-EVAL: endmodule not found
