
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
localparam B = 1'b1;
localparam A = 1'b0;

reg state, next_state;

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= B;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        B: next_state = in ? B : A;
        A: next_state = in ? A : B;
        default: next_state = B;
    endcase
end

assign out = state;

endmodule
