
module TopModule (
  input cpu_overheated,
  output reg shut_off_computer,
  input arrived,
  input gas_tank_empty,
  output reg keep_driving
);
module top_module (
    input cpu_overheated,
    output reg shut_off_computer,
    input arrived,
    input gas_tank_empty,
    output reg keep_driving
);

always @(posedge clk) begin // Added posedge clause for proper synchronization
    if (cpu_overheated)
        shut_off_computer <= 1;
end

always @(posedge clk) begin // Added posedge clause for proper synchronization
    if (!arrived)
        keep_driving <= !gas_tank_empty;
end

endmodule
