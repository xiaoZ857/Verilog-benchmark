
module TopModule (
  input a,
  input b,
  input c,
  output w,
  output x,
  output y,
  output z
);


// VERILOG-EVAL: endmodule not found
