

module TopModule (
  input clk,
  input reset,
  output [3:1] ena,
  output reg [15:0] q
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        q <= 16'b0000_0000_0000_0000;
        ena <= 3'b000;
    end else begin
        // Increment the ones digit
        if (q[3:0] == 4'd9) begin
            q[3:0] <= 4'd0;
            ena[1] <= 1'b1; // Enable tens digit increment
        end else begin
            q[3:0] <= q[3:0] + 1;
            ena[1] <= 1'b0;
        end

        // Increment the tens digit
        if (q[7:4] == 4'd9) begin
            q[7:4] <= 4'd0;
            ena[2] <= 1'b1; // Enable hundreds digit increment
        end else if (ena[1]) begin
            q[7:4] <= q[7:4] + 1;
            ena[2] <= 1'b0;
        end

        // Increment the hundreds digit
        if (q[11:8] == 4'd9) begin
            q[11:8] <= 4'd0;
            ena[3] <= 1'b1; // Enable thousands digit increment
        end else if (ena[2]) begin
            q[11:8] <= q[11:8] + 1;
            ena[3] <= 1'b0;
        end

        // Increment the thousands digit
        if (ena[3]) begin
            if (q[15:12] == 4'd9) begin
                q[15:12] <= 4'd0; // Reset to zero after reaching 9999
            end else begin
                q[15:12] <= q[15:12] + 1;
            end
        end
    end
end

// Ensure ena is always driven correctly
always @(*) begin
    if (q[3:0] == 4'd9) ena[1] = 1'b1;
    else ena[1] = 1'b0;

    if (q[7:4] == 4'd9) ena[2] = 1'b1;
    else ena[2] = 1'b0;

    if (q[11:8] == 4'd9) ena[3] = 1'b1;
    else ena[3] = 1'b0;
end

endmodule
