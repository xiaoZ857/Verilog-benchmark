
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);
reg [1:0] state;
reg [1:0] next_state;

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= 2'b01; // Reset to state A
    else
        state <= next_state;
end

always @* begin
    case (state)
        2'b01: // State A
            next_state = x ? 2'b10 : 2'b01;
        2'b10: // State B
            next_state = 2'b10;
        default:
            next_state = 2'b01;
    endcase
end

assign z = state[0] ? x : ~x;

endmodule
