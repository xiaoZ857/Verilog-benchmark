
module TopModule (
  input a,
  input b,
  input c,
  output out
);
out = a | b | c;

// VERILOG-EVAL: endmodule not found
