
  always @(*) begin
      case (do_sub)
        0: out = a+b;
        1: out = a-b;
      endcase

      if (out == 8'b0)
          result_is_zero = 1;
      else
          result_is_zero = 0;
  end

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
