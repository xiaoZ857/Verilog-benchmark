

module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);



// VERILOG-EVAL: endmodule not found
