
// Assign 0 to the output 'zero' continuously
assign zero = 0;

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
