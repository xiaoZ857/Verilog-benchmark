
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  output walk_left,
  output walk_right,
  output aaah
);

reg [1:0] state, next_state;

// State encoding
parameter WALK_LEFT  = 2'b00;
parameter WALK_RIGHT = 2'b01;
parameter FALL_LEFT  = 2'b10;
parameter FALL_RIGHT = 2'b11;

// State register
always @(posedge clk or posedge areset) begin
    if (areset)
        state <= WALK_LEFT;
    else
        state <= next_state;
end

// Next state logic
always @(*) begin
    case (state)
        WALK_LEFT: begin
            if (ground == 0)
                next_state = FALL_LEFT;
            else if (bump_left)
                next_state = WALK_RIGHT;
            else
                next_state = WALK_LEFT;
        end
        
        WALK_RIGHT: begin
            if (ground == 0)
                next_state = FALL_RIGHT;
            else if (bump_right)
                next_state = WALK_LEFT;
            else
                next_state = WALK_RIGHT;
        end
        
        FALL_LEFT: begin
            if (ground == 1)
                next_state = WALK_LEFT;
            else
                next_state = FALL_LEFT;
        end
        
        FALL_RIGHT: begin
            if (ground == 1)
                next_state = WALK_RIGHT;
            else
                next_state = FALL_RIGHT;
        end
        
        default: next_state = WALK_LEFT;
    endcase
end

// Output logic (Moore machine - outputs depend only on state)
assign walk_left  = (state == WALK_LEFT);
assign walk_right = (state == WALK_RIGHT);
assign aaah = (state == FALL_LEFT) || (state == FALL_RIGHT);

endmodule
