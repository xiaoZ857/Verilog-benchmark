
module TopModule (
  input wire in,
  output wire out
);

  // Combinational assignment of the output to the input
  assign out = in;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
