

module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);

  // State encoding
  // 3'd0 : SEARCH  �C look for a byte with in[3]==1
  // 3'd

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
