
module TopModule (
  input clk,
  input reset,
  output reg [9:0] q
);
always @(posedge clk or posedge reset) begin
    if (reset)
        q <= 10'd0;
    else
        q <= (q == 10'd999) ? 10'd0 : q + 1'b1;
end
endmodule
