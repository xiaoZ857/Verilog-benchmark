
module TopModule (
  input in,
  output out
);
  
  // Assign input 'in' directly to output 'out'
  assign out = in;
  
endmodule

// VERILOG-EVAL: errant inclusion of module definition
