
module TopModule (
  input [1023:0] in,
  input [7:0] sel,
  output [3:0] out
);
  out = in[sel*4 +: 4];

// VERILOG-EVAL: endmodule not found
