
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);

  // State encoding
  parameter A = 3'b000;
  parameter B = 3'b001;
  parameter C = 3'b010;
  parameter D = 3'b011;
  parameter E = 3'b100;
  parameter F = 3'b101;
  
  // State registers
  reg [2

// VERILOG-EVAL: endmodule not found
