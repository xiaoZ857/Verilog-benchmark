
module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);
always @(posedge clk or posedge reset) // Combining both positive edges for clock and reset
begin
    if (reset) begin
        q <= 4'b0001; // Reset value is 1 (decimal 1, binary 0001)
    end else begin
        if (q == 4'b1001) begin // Check if counter reaches the maximum value of 10 (decimal)
            q <= 4'b0001; // Reset counter to start counting again
        end else begin
            q <= {q[3], q[2]+1'b0, q[1], q[0]+1'b0}; // Shift left and increment lower bits (casting q[2] and q[0] to 1-bit)
        end
    end
end

// Testbench for TopModule verification
module testbench;

reg clk, reset;
wire [3:0] q;
TopModule uut (clk, reset, q);

initial begin
    always #5 clk = ~clk; // Generate a clock signal with 5ns period

    // Initialization
    reset = 0;
    #10;
    reset = 1; // Reset the counter at time 10ns

    // Simulation for 60ns to observe counter behavior
    #40 $finish;
end

// VERILOG-EVAL: endmodule not found
