
module TopModule (
  input [7:0] in,
  output [7:0] out
);

assign out[0] = in[7];
assign out[1] = in[6];
assign

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
