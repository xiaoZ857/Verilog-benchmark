
// 10‑state decade counter (0 … 9)
//  - synchronous active‑high reset
//  - "slowena" enables increment on each clock edge
module TopModule (
    input  wire        clk,      // clock
    input  wire        slowena,  // enable increment
    input  wire        reset,    // active‑high synchronous reset
    output reg  [3:0]  q         // 4‑bit counter output
);

    // synchronous logic
    always @(posedge clk) begin
        if (reset) begin
            // synchronous reset – takes priority over slowena
            q <= 4'd0;
        end
        else if (slowena) begin
            // increment only when enabled
            if (q == 4'd9) begin
                q <= 4'd0;        // wrap‑around
            end else begin
                q <= q + 1'b1;    // normal increment
            end
        end
        // else: retain current value (paused)
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
