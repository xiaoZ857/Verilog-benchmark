
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
  reg state;
  localparam B = 1'b0, A = 1'b1;
  
  always @(posedge clk) begin
    if (reset) begin
      state <= B;
    end else begin
      case (state)
        B: state <= in ? B : A;
        A: state <= in ? A : B;
        default: state <= B;
      endcase
    end
  end
  
  assign out = (state == B) ? 1'b1 : 1'b0;
endmodule
