
module TopModule (
  input clk,
  input enable,
  input S,
  input A,
  input B,
  input C,
  output reg Z
);
always @(posedge clk) begin
    if (enable) begin
        Z <= {Z[6:0], S};
    end
end

always @(*) begin
    case ({A, B, C})
        3'b000: Z = Z[0];
        3'b001: Z = Z[1];
        3'b010: Z = Z[2];
        3'b011: Z = Z[3];
        3'b100: Z = Z[4];
        3'b101: Z = Z[5];
        3'b110: Z = Z[6];
        3'b111: Z = Z[7];
        default: Z = 1'b0;
    end
end

endmodule
