

module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);

reg [1:0] current_state, next_state;

localparam S0 = 2'b00;
localparam S1 = 2'b01;
localparam S2 = 2'b10;

always @(posedge clk or negedge aresetn) begin
    if (!aresetn)
        current_state <= S0;
    else
        current_state <= next_state;
end

always @(*) begin
    case (current_state)
        S0: 
            if (x == 1'b1)
                next_state = S1;
            else
                next_state = S0;

        S1:
            if (x == 1'b0)
                next_state = S2;
            else
                next_state = S1;

        S2:
            if (x == 1'b1)
                next_state = S1;
            else
                next_state = S0;

        default: 
            next_state = S0;
    endcase
end

always @(posedge clk or negedge aresetn) begin
    if (!aresetn)
        z <= 1'b0;
    else begin
        case (current_state)
            S2:
                if (x == 1'b1)
                    z <= 1'b1;
                else
                    z <= 1'b0;

            default: 
                z <= 1'b0;
        endcase
    end
end

endmodule
