

module TopModule (
  input x,
  input y,
  output z
);

assign z = (x'1 && ~y) || (~x & y);
endmodule
