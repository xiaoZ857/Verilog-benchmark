

module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);



// VERILOG-EVAL: endmodule not found
