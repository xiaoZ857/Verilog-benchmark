
module TopModule (
  input [15:0] scancode,
  output reg left,
  output reg down,
  output reg right,
  output reg up
);

  always @(scancode) begin
    left = 0;
    down = 0;
    right = 0;
    up = 0;

    case (scancode)
      16'h06b: left = 1;
      16'h072: down = 1;
      16'h074: right = 1;
      16'h075: up = 1;
      default: ; // Do nothing if not an arrow key
    endcase
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
