
module TopModule (
    input  wire        clk,        // clock
    input  wire        shift_ena,  // shift enable
    input  wire        count_ena,  // count enable
    input  wire        data,       // data to shift in (MSB first)
    output reg  [3:0]  q           // 4‑bit register
);

    // S

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
