

module TopModule (
  input a,
  input b,
  output q
);

  always @(a or b) begin
    if (a == 0 && b == 0) begin
      q = 0;
    end else if (a == 0 && b == 1) begin
      q = 0;
    end else if (a == 1 && b == 0) begin
      q = 0;
    end else begin
      q = 1;
    end
  end
endmodule
