

module TopModule (
  input [255:0] in,
  input [7:0] sel,
  output  out
);

always @(posedge clk) begin
    case (sel)
        8'b00000000: out <= in[0];
        8'b00000001: out <= in[1];
        8'b00000010: out <= in[2];
        8'b00000011: out <= in[3];
        8'b00000100: out <= in[4];
        8'b00000101: out <= in[5];
        8'b00000110: out <= in[6];
        8'b00000111: out <= in[7];
        8'b00001000: out <= in[8];
        8'b00001001: out <= in[9];
        8'b00001010: out <= in[10];
        8'b00001011: out <= in[11];
        8'b00001100: out <= in[12];
        8'b00001101: out <= in[13];
        8'b00001110: out <= in[14];
        8'b00001111: out <= in[15];
        8'b00010000: out <= in[16];
        8'b00010001: out <= in[17];
        8'b00010010: out <= in[18];
        8'b00010011: out <= in[19];
        8'b00010100: out <= in[20];
        8'b00010101: out <= in[21];
        8'b00010110: out <= in[22];
        8'b00010111: out <= in[23];
        8'b00011000: out <= in[24];
        8'b00011001: out <= in[25];
        8'b00011010: out <= in[26];
        8'b00011011: out <= in[27];
        8'b00011100: out <= in[28];
        8'b00011101: out <= in[29];
        8'b00011110: out <= in[30];
        8'b00011111: out <= in[31];
        8'b00100000: out <= in[32];
        8'b00100001: out <= in[33];
        8'b00100010: out <= in[34];
        8'b00100011: out <= in[35];
        8'b00100100: out <= in[36];
        8'b00100101: out <= in[37];
        8'b00100110: out <= in[38];
        8'b00100111: out <= in[39];
        8'b00101000: out <= in[40];
        8'b00101001: out <= in[41];
        8'b00101010: out <= in[42];
        8'b00101011: out <= in[43];
        8'b00101100: out <= in[44];
        8'b00101101: out <= in[45];
        8'b00101110: out <= in[46];
        8'b00101111: out <= in[47];
        8'b00110000: out <= in[48];
        8'b00110001: out <= in[49];
        8'b00110010: out <= in[50];
        8'b00110011: out <= in[51];
        8'b00110100: out <= in[52];
        8'b00110101: out <= in[53];
        8'b00110110: out <= in[54];
        8'b00110111: out <= in[55];
        8'b00111000: out <= in[56];
        8'b00111001: out <= in[57];
        8'b00111010: out <= in[58];
        8'b00111011: out <= in[59];
        8'b00111100: out <= in[60];
        8'b00111101: out <= in[61];
        8'b00111110: out <= in[62];
        8'b00111111: out <= in[63];
        8'b01000000: out <= in[64];
        8'b01000001: out <= in[65];
        8'b01000010: out <= in[66];
        8'b01000011: out <= in[67];
        8'b01000100: out <= in[68];
        8'b01000101: out <= in[69];
        8'b01000110: out <= in[70];
        8'b01000111: out <= in[71

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
