
      ab
   cd  00  01  11  10
   00 | 1 | 1 | 0 | 1 |
   01 | 1 | 0 | 0 | 1 |
   11 | 0 | 1 | 1 | 1 |
   10 | 1 | 1 | 0 | 0 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
