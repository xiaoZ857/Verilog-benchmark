
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);
// Define the states of the Lemming FSM
parameter [1:0] stateWalking = 2'b00;
parameter [1:0] stateDigging = 2'b01;
parameter [1:0] stateFalling = 2'b10;

// Define the next state for each input transition
localparam NEXT_STATE_WALKING_BUMP_LEFT = stateWalking + 1'b1;
localparam NEXT_STATE_DIGGING_BUMP_LEFT = stateWalking; 
localparam NEXT_STATE_FALLING_BUMP_LEFT = stateFalling;

localparam NEXT_STATE_WALKING_BUMP_RIGHT = stateWalking - 1'b1;
localparam NEXT_STATE_DIGGING_BUMP_RIGHT = stateWalking; 
localparam NEXT_STATE_FALLING_BUMP_RIGHT = stateFalling;

// Define the state machines for falling and digging
parameter [2:0] FALLING_STATE = 3'b100;
parameter [2:0] DIGGING_STATE = 3'b000;

parameter [2:0] NEXT_FALLING_STATE = {stateFalling, fallCounter};
parameter [2:0] NEXT_DIGGING_STATE = {stateDigging, digCounter};

// Initialize counters for falling and digging
wire [1:0] fallCounter;
wire [1:0] digCounter;

assign fallCounter = ~falling_state[2'b00];

// Initialize digging state machine with a counter
RegNext stateDiggingReg(\~dig);
RegNext nextStateDiggingReg(\stateDigging);

assign nextStateDiggingReg.NEXT_STATE = NEXT_DIGGING_STATE;
assign stateDiggingReg.NEXT_STATE = NEXT_STATE DIGGING_BUMP_LEFT; // Corrected to only bump left

// Initialize falling state machine with a counter
RegNext stateFallingReg(\~ground);
RegNext nextStateFallingReg(\stateFalling);

assign nextStateFallingReg.NEXT_STATE = NEXT_FALLING_STATE;
assign stateFallingReg.NEXT_STATE = NEXT_STATE_FALLING_BUMP_LEFT; // Corrected to only bump left

// Initialize walk_left and walk_right outputs
wire walkLeftOutput;
wire walkRightOutput;

RegNext nextStateWalkingReg(\stateWalking);
RegNext nextNextStateWalkingReg(NEXT_STATE_WALKING_BUMP_LEFT, NEXT_STATE_WALKING_BUMP_RIGHT, NEXT_STATE_FALLING_BUMP_LEFT);

assign nextNextStateWalkingReg.NEXT_STATE = nextStateWalkingReg.NEXT_STATE;
assign walkLeftOutput = (nextNextStateWalkingReg == stateWalking + 1'b1) ? 1'b0 : (nextNextStateWalkingReg == stateWalking - 1'b1) ? 1'b1 : 0'b0;

// Initialize aaah output
RegNext nextStateAAahReg(\~ground);
RegNext nextNextStateAAahReg(NEXT_STATE_FALLING);

assign nextNextStateAAahReg.NEXT_STATE = nextStateAAahReg.NEXT_STATE;
assign aaah = (nextNextStateAAahReg == stateWalking) ? 1'b0 : 1'b1;

// Asynchronous reset
RegNext nextStateAAahReg_AsyncReset(NEXT_STATE_FALLING);

RegNext nextStateWalkingDigReg_NextState(\~dig);
RegNext nextStateWalkingDigRegNEXT_STATE(NEXT_STATE_WALKING_BUMP_LEFT, NEXT_STATE_WALKING_BUMP_RIGHT, NEXT_STATE_FALLING_BUMP_LEFT);

assign nextStateWalkingDigRegNEXT_STATE.NEXT_STATE = nextStateWalkingDigReg.NEXT_STATE;
assign walkRightOutput = (nextStateWalkingDigRegNEXT_STATE == stateWalking - 1'b1) ? 1'b0 : 0'b0;

// Assignments for digging
RegNext nextStateDiggingReg (\stateDigging);
RegNext nextNextStateDiggingReg(NEXT_STATE_DIGGING_BUMP_LEFT, NEXT_STATE_DIGGING_BUMP_RIGHT, NEXT_STATE_FALLING_BUMP_LEFT);

assign nextStateDiggingReg.NEXT_STATE = nextNextStateDiggingReg.NEXT_STATE;

// Asynchronous reset for digging
RegNext digResetReg (\~reset);
RegNext nextStateDiggingReg_NextState_Digreset(\~dig, \reset);

assign nextStateDiggingReg_NextState_Digreset.NEXT_STATE = nextStateDiggingReg.NEXT_STATE;
assign digResetReg.NEXT_STATE = NEXT_STATE_DIGGING_BUMP_LEFT;

// Counters for digging
wire [1:0] digCounter;

assign digCounter = ~digResetReg;

// Splatter detection
wire splatter;
assign splatter = fallCounter[2'b00] == 20'b000 && stateWalkingReg.NEXT_STATE == stateFallingReg.NEXT_STATE;

// Reset FSM when Lemming splatters or falls for too long
RegNext nextStateLemmingReg(\~splatter);
RegNext nextStateAAahReg(\~splatter);
RegNext nextNextStateLemmingReg(NEXT_STATE_FALLING, NEXT_STATE SPLATTERED);

assign nextNextStateLemmingReg.NEXT_STATE = nextStateLem

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
