
module TopModule (
  input [99:0] in,
  output [98:0] out_both,
  output [99:1] out_any,
  output [99:0] out_different
);
always_comb begin
    // Calculate out_both
    for (int i = 0; i < 98; i++) begin
        out_both[i] = in[i] & in[i + 1];
    end

    // Calculate out_any
    for (int i = 2; i <= 99; i++) begin
        out_any[i - 2] = in[i - 1] | in[i];
    end

    // Calculate out_different
    for (int i = 0; i < 100; i++) begin
        int left_index = (i + 1) % 100;
        out_different[i] = in[i] != in[left_index];
    end
endmodule

// VERILOG-EVAL: abnormal backticks count
