
module TopModule(
    input clk,            // Positive edge triggered clock signal
    input [7:0] in,         // Byte stream with MSB on top
    input reset,           // Asynchronous active high reset signal
    output done             // Signal indicating message has been received
);

// Internal signals for the state machine
reg [2:0] state;
reg [7:0] messageBytes[3];  // Storing the last 3 bytes of a message

// Constructor for the state machine
always @(posedge clk or negedge reset) begin
    if(reset)
        state <= 2;      // Reset to idle state
    else
        case(state)
            0: state <= 1;    // Start byte detected, start searching for message boundary
            1: state <= 2;
            2: state <= 3;    // Message boundary found, start reading the first byte of a message
            3: state <= 0;    // First byte of a message read, start reading the second byte
            default: state <= 0;
        endcase
end

// Reading bytes from the input stream and checking if they form a valid message
always @(posedge clk or (in[7] == 1)) begin
    if(state == 3) begin
        if(in[7:0] == messageBytes[2])   // Check if second byte matches the last one of the previous message
            state <= 4;                  // Continue reading the third and final byte of a message
        else
            state <= 0;
    end
    else if(state == 4) begin
        if(in[7:0] == messageBytes[3])   // Check if last one of this message matches the second to last of previous one's (message boundary)
            done <= 1;                   // A full message has been received
        else
            state <= 0;
    end
end

// Writing the bytes to internal memory and signaling when a message is read
always @(posedge clk) begin
    if(state == 4) begin
        messageBytes[3] <= in[7:0];
        done <= 1;
    end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
