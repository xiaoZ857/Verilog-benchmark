

module TopModule (
  input clk,
  input reset,
  output reg [9:0] q
);



// VERILOG-EVAL: endmodule not found
