
module TopModule (
  output out
);
  assign out = 1'b0;
endmodule

// VERILOG-EVAL: errant inclusion of module definition
