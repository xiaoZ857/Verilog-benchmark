
// TopModule.v
// 7‑output combinational logic – each output is produced by a single logic gate.

module TopModule (
    input  wire a,          // first input
    input  wire b,          // second input
    output wire out_and,    // a AND b
    output wire out_or,     // a OR  b
    output wire out_xor,    // a XOR b
    output wire out_nand,   // a NAND b
    output wire out_nor,    // a NOR  b
    output wire out_xnor,   // a XNOR b
    output wire out_anotb   // a AND NOT b
);

    // ----- Gate instantiations ---------------------------------
    and  g_and    (out_and,  a, b);           // a & b
    or   g_or     (out_or,   a, b);           // a | b
    xor  g_xor    (out_xor,  a, b);           // a ^ b
    nand g_nand   (out_nand, a, b);           // ~(a & b)
    nor  g_nor    (out_nor,  a, b);           // ~(a | b)
    xnor g_xnor   (out_xnor, a, b);           // ~(a ^ b)
    and  g_anotb  (out_anotb, a, ~b);         // a & (~b)

    // (Optional) you could also write the same logic with continuous assignments:
    // assign out_and   = a & b;
    // assign out_or    = a | b;
    // assign out_xor   = a ^ b;
    // assign out_nand  = ~(a & b);
    // assign out_nor   = ~(a | b);
    // assign out_xnor  = ~(a ^ b);
    // assign out_anotb = a & ~b;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
