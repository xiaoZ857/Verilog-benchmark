
module TopModule (
    input wire clk,
    input wire [7:0] in,
    input wire reset,
    output reg [23:0] out_bytes,
    output reg done
);

    // State encoding
    typedef enum logic [1:0] {
        IDLE = 2'b00,  // Waiting for start byte
        RECV_BYTE_1 = 2'b01,  // Receiving first byte of message
        RECV_BYTE_2 = 2'b10,  // Receiving second byte of message
        RECV_BYTE_3 = 2'b11   // Receiving third byte of message
    } state_t;

    state_t current_state, next_state;
    
    reg [7:0] byte1, byte2;  // Registers to store the first two bytes

    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            current_state <= IDLE;
            done <= 0;
            out_bytes <= 24'b0;
        end else begin
            current_state <= next_state;

            case (current_state)
                RECV_BYTE_1: begin
                    byte1 <= in;
                end
                RECV_BYTE_2: begin
                    byte2 <= in;
                end
                RECV_BYTE_3: begin
                    out_bytes <= {byte1, byte2, in};
                    done <= 1;
                end
            endcase

            // Reset the 'done' signal only after the output has been latched
            if (current_state == RECV_BYTE_3) begin
                done <= 0;
            end
        end
    end

    always_comb begin
        next_state = current_state;  // Default to stay in same state
        case (current_state)
            IDLE: begin
                if (in[3]) begin
                    next_state = RECV_BYTE_1;
                end
            end
            RECV_BYTE_1: begin
                next_state = RECV_BYTE_2;
            end
            RECV_BYTE_2: begin
                next_state = RECV_BYTE_3;
            end
            RECV_BYTE_3: begin
                next_state = IDLE;  // Return to idle after receiving a message
            end
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
