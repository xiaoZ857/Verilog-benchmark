
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out
);
    // Always block to be triggered on each clock edge
    always @(posedge clk) begin
        // Karnaugh map implementation:
        // ab  cd   00  01  11  10
        // 00 | 1 | 1 | 0 | 1 |
        // 01 | 1 | 0 | 0 | 1 |
        // 11 | 0 | 1 | 1 | 1 |
        // 10 | 1 | 1 | 0 | 0 |

        out <= (a & b) | ((c & d) | (~c & ~d)); // Applying De Morgan's laws
    end
endmodule
