
module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);
always @(posedge clk or negedge aresetn) begin
    if (!aresetn) begin
        z <= 1'b0;
    end else begin
        case (state)
            S0: begin
                if (x) begin
                    state <= S1;
                    z <= 1'b0;
                end else begin
                    state <= S0;
                    z <= 1'b0;
                end
            end
            S1: begin
                if (!x) begin
                    state <= S2;
                    z <= 1'b0;
                end else begin
                    state <= S1;
                    z <= 1'b0;
                end
            end
            S2: begin
                if (x) begin
                    state <= S1;
                    z <= 1'b1;
                end else begin
                    state <= S0;
                    z <= 1'b0;
                end
            end
            default: begin
                state <= S0;
                z <= 1'b0;
            end
        endcase
    end
end

reg [1:0] state;
parameter S0 = 2'b00, S1 = 2'b01, S2 = 2'b10;

endmodule
