
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
reg [1:0] state, next_state;

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= 2'b00; // Reset to state A
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        2'b00: begin // State A
            out = 1'b0;
            if (in == 1'b0) 
                next_state = 2'b00; // Remain in state A
            else
                next_state = 2'b01; // Transition to state B
        end
        2'b01: begin // State B
            out = 1'b0;
            if (in == 1'b0)
                next_state = 2'b10; // Transition to state C
            else
                next_state = 2'b01; // Remain in state B
        end
        2'b10: begin // State C
            out = 1'b0;
            if (in == 1'b0)
                next_state = 2'b00; // Transition to state A
            else
                next_state = 2'b11; // Transition to state D
        end
        2'b11: begin // State D
            out = 1'b1;
            if (in == 1'b0)
                next_state = 2'b10; // Transition to state C
            else
                next_state = 2'b01; // Transition to state B
        end
    endcase
end

endmodule
