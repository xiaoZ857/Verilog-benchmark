
module TopModule (
  input p1a,
  input p1b,
  input p1c,
  input p1d,
  output p1y,
  input p2a,
  input p2b,
  input p2c,
  input p2d,
  output p2y
);

  // NAND gate 1: p1y = NOT(p1a AND p1b AND p1c AND p1d)
  assign p1y = ~ (p1a & p1b & p1c & p1d);

  // NAND gate 2: p2y = NOT(p2a AND p2b AND p2c AND p2d)
  assign p2y = ~ (p2a & p2b & p2c & p2d);

endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
