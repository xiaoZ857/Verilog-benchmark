

module TopModule (
  input clk,
  input d,
  output reg q
);

always @(posedge clk) begin
  if (d) begin
    q <= 1;
  end else begin
    q <= 0;
  end
end

always @(negedge clk) begin
  if (d) begin
    q <= 1;
  end else begin
    q <= 0;
  end
end

endmodule
