
module TopModule (
  input clk,
  input areset,
  input train_valid,
  input train_taken,
  output logic [1:0] state
);
always @(posedge clk) begin
    if (areset) begin
        state <= 2'b01; // Asynchronous reset sets counter to weakly not-taken (2'b01)
    end else if (train_valid && train_taken) begin
        state <= state + 1; // Increment counter up to maximum of 3
        if (state > 3'b11) state <= 3'b11; // Saturating at maximum value
    end else if (train_valid && !train_taken) begin
        state <= state - 1; // Decrement counter down to minimum of 0
        if (state < 2'b00) state <= 2'b00; // Saturating at minimum value
    end
end

// Adding timescale directive outside the module definition as requested.
`timescale 1ns / 1ps

// VERILOG-EVAL: endmodule not found
