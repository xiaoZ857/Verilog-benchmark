
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output reg out
);
out = a'b'c + a'bcd'

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
