
//  Two‑bit saturating counter
//  state  : 2‑bit value (00 … 11)
//  areset : asynchronous reset (active‑high)
//  clk    : synchronous clock
//  train_valid : enable for training
//  train_taken : direction of the update
//
//  Behaviour
//    • If areset is asserted – state is reset to 2'b01 (weakly “not‑taken”).
//    • When train_valid = 1
//          – if train_taken = 1 : increment (saturate at 3)
//          – if train_taken = 0 : decrement (saturate at 0)
//    • When train_valid = 0 : keep the current state.

module TopModule (
    input  logic        clk,
    input  logic        areset,
    input  logic        train_valid,
    input  logic        train_taken,
    output logic [1:0]  state
);

    // The counter is updated on the rising edge of clk.
    // The asynchronous reset is also taken into account.
    always_ff @(posedge clk or posedge areset)
    begin
        if (areset) begin
            // Asynchronous reset – initialise to weakly not‑taken
            state <= 2'b01;
        end
        else if (train_valid) begin
            // Only update when training is active
            if (train_taken) begin
                // Increment but saturate at 3 (binary 11)
                if (state != 2'b11)
                    state <= state + 1'b1;
            end
            else begin
                // Decrement but saturate at 0 (binary 00)
                if (state != 2'b00)
                    state <= state - 1'b1;
            end
        end
        // If train_valid == 0 → state stays unchanged
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
