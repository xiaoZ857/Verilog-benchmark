

module TopModule (
  input clk,
  input load,
  input [9:0] data,
  output tc
);



// VERILOG-EVAL: endmodule not found
