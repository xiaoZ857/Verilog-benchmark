
      even number of 1’s  →  q = 1
      odd  number of 1’s  →  q = 0

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
