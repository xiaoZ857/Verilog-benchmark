

module TopModule (
  input [2:0] sel,
  input [3:0] data0,
  input [3:0] data1,
  input [3:0] data2,
  input [3:0] data3,
  input [3:0] data4,
  input [3:0] data5,
  output reg [3:0] out
);

always @(posedge clk) begin
  case (sel)
    2'b00 : out <= data0;
    2'b01 : out <= data1;
    2'b10 : out <= data2;
    2'b110 : out <= data3;
    2'b1110 : out <= data4;
    2'b11110 : out <= data5;
    default : out <= 4'b0000; // Output 0 when sel is not between 0 and 5
  endcase
end

// VERILOG-EVAL: endmodule not found
