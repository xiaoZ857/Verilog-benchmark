
module TopModule (
    input  wire        in,          // asynchronous input
    input  wire [3:0]  state,       //

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
