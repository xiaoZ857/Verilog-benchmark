

module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

reg [2:0] state, next_state;

localparam IDLE_LEFT = 3'b000;
localparam WALK_RIGHT = 3'b001;
localparam FALLING = 3'b010;
localparam DIGGING = 3'b011;
localparam IDLE_RIGHT = 3'b100;

assign walk_left = (state == IDLE_LEFT) | (state == FALLING) | (state == DIGGING);
assign walk_right = (state == WALK_RIGHT) | (state == IDLE_RIGHT) | (state == FALLING) | (state == DIGGING);
assign aaah = (state == FALLING) | (state == DIGGING);
assign digging = (state == DIGGING);

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= IDLE_LEFT;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        IDLE_LEFT: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_left || bump_right)
                next_state = WALK_RIGHT;
            else if (dig)
                next_state = DIGGING;
            else
                next_state = IDLE_LEFT;
        end

        WALK_RIGHT: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_left || bump_right)
                next_state = IDLE_LEFT;
            else
                next_state = WALK_RIGHT;
        end

        FALLING: begin
            if (ground)
                next_state = state == IDLE_LEFT ? IDLE_LEFT : IDLE_RIGHT;
            else
                next_state = FALLING;
        end

        DIGGING: begin
            if (!ground)
                next_state = FALLING;
            else if (ground && !dig)
                next_state = state == IDLE_LEFT ? IDLE_LEFT : IDLE_RIGHT;
            else
                next_state = DIGGING;
        end

        IDLE_RIGHT: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_left || bump_right)
                next_state = WALK_LEFT;
            else if (dig)
                next_state = DIGGING;
            else
                next_state = IDLE_RIGHT;
        end

        default: next_state = IDLE_LEFT;
    endcase
end

endmodule
