
module TopModule (
  input [7:0] code,
  output reg [3:0] out,
  output reg valid
);


// VERILOG-EVAL: endmodule not found
