
module TopModule (
    input  wire clk,   // positive‑edge clock
    input  wire x,     // data input
    output wire z      // FSM output
);

    // Flip‑flop outputs (state)
    reg q0, q1, q2;

    // Initialise the state to 0 (

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
