
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);


// VERILOG-EVAL: endmodule not found
