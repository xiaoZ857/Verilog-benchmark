
module TopModule (
  output one
);
assign one = 1;

// VERILOG-EVAL: endmodule not found
