
module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);
always @(posedge clk) begin
    if (load) begin
        q <= data;
    end else begin
        
        logic [255:0] next_q;
        
        for (int i = 0; i < 256; i++) begin
            logic neighbors;
            
            // Get the current cell value
            logic current_cell = q[i];
            
            // Calculate the number of neighbors
            neighbors = 0;
            
            // Wrap-around logic for neighbor calculation
            for (int j = -1; j <= 1; j++) {
                for (int k = -1; k <= 1; k++) {
                    if (j == 0 && k == 0) continue;
                    
                    int neighbor_index = i + j * 16 + k;
                    
                    if (neighbor_index < 0) neighbor_index += 256;
                    if (neighbor_index >= 256) neighbor_index -= 256;
                    
                    neighbors = neighbors | q[neighbor_index];
                }
            }
            
            // Update the cell based on the game rules
            if (neighbors == 1)
                next_q[i] = 0;
            else if (neighbors == 2)
                next_q[i] = current_cell;
            else if (neighbors == 3)
                next_q[i] = 1;
            else if (neighbors >= 4)
                next_q[i] = 0;
            else
                next_q[i] = current_cell;
        }
        q <= next_q;
    end
endmodule
