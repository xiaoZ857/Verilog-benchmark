
module TopModule (
  input clk,
  input reset,
  input data,
  output reg shift_ena,
  output reg counting,
  input done_counting,
  output reg done,
  input ack
);

  // State encoding
  typedef enum logic [2:0] {
    IDLE       = 3'b000,  // Waiting for start sequence
    DETECT_1   = 3'b001,  // Detected '1' in sequence
    DETECT_11  = 3'b010,  // Detected '11' in sequence
    DETECT_110 = 3'b011,  // Detected '110' in sequence
    START      = 3'b100,  // Detected start pattern '1101'
    SHIFT      = 3'b101,  // Shifting the next 4 bits for delay
    COUNT      = 3'b110,  // Waiting for counters to finish
    NOTIFY     = 3'b111   // Notifying user and waiting for acknowledgment
  } state_t;

  state_t current_state, next_state;

  always_ff @(posedge clk or posedge reset) begin
    if (reset)
      current_state <= IDLE;
    else
      current_state <= next_state;
  end

  always_comb begin
    // Default outputs and next state
    shift_ena = 1'b0;
    counting = 1'b0;
    done = 1'b0;
    next_state = current_state;

    case (current_state)
      IDLE: begin
        if (data == 1'b1) 
          next_state = DETECT_1;
      end

      DETECT_1: begin
        if (data == 1'b1)
          next_state = DETECT_11;
        else
          next_state = IDLE;
      end

      DETECT_11: begin
        if (data == 1'b0)
          next_state = DETECT_110;
        else
          next_state = DETECT_1;
      end

      DETECT_110: begin
        if (data == 1'b1)
          next_state = START;
        else
          next_state = IDLE;
      end

      START: begin
        shift_ena = 1'b1; // Enable shifting of the next 4 bits
        next_state = SHIFT;
      end

      SHIFT: begin
        shift_ena = 1'b0; // Disable shifting after 4 cycles
        if (data) 
          next_state = COUNT; // Shifted all 4 bits, proceed to counting
      end

      COUNT: begin
        counting = 1'b1; // Start counting
        if (done_counting)
          next_state = NOTIFY;
      end

      NOTIFY: begin
        done = 1'b1; // Notify the user
        if (ack)
          next_state = IDLE; // Wait for acknowledgment and reset
      end
      
    endcase
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
