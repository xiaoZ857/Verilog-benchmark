
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  output walk_left,
  output walk_right
);
// State encoding for the two possible states
parameter WALK_LEFT = 1'b0;
parameter WALK_RIGHT = 1'b1;

reg current_state;
reg next_state;

// State transition logic
always @(*) begin
  case (current_state)
    WALK_LEFT: begin
      if (bump_left) begin
        next_state = WALK_RIGHT;
      end else begin
        next_state = WALK_LEFT;
      end
    end
    WALK_RIGHT: begin
      if (bump_right) begin
        next_state = WALK_LEFT;
      end else begin
        next_state = WALK_RIGHT;
      end
    end
    default: next_state = WALK_LEFT;
  endcase
end

// State update and reset logic
always @(posedge clk or posedge areset) begin
  if (areset) begin
    current_state <= WALK_LEFT;
  end else begin
    current_state <= next_state;
  end
end

// Output logic (Moore machine - outputs depend only on current state)
assign walk_left = (current_state == WALK_LEFT);
assign walk_right = (current_state == WALK_RIGHT);

endmodule
