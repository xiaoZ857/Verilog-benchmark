
module TopModule (
  input a,
  input b,
  output q
);

// Implementing the AND function
q = a & b;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
