
module TopModule (
  input clk,
  input a,
  input b,
  output out_assign,
  output reg out_always_comb,
  output reg out_always_ff
);

  // Implement XOR using an assign statement (combinational logic)
  assign out_assign = a ^ b;

  // Implement XOR using a combinational always block
  always @(*) begin
    out_always_comb = a ^ b;
  end

  // Implement XOR using a clocked always block with a flip-flop
  always @(posedge clk) begin
    out_always_ff <= a ^ b;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
