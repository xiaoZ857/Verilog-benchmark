
module TopModule (
    input [4:0] a,
    input [4:0] b,
    input [4:0] c,
    input [4:0] d,
    input [4:0] e,
    input [4:0] f,
    output [7:0] w,
    output [7:0] x,
    output [7:0] y,
    output [7:0] z
);

    // Concatenate the input vectors into a 30-bit vector
    wire [29:0] inputVector = {a, b, c, d, e, f};

    // Split the input vector into four 8-bit vectors
    assign w[7:0] = inputVector[24:15];
    assign x[7:0] = inputVector[20:11];
    assign y[7:0] = inputVector[16:7];
    assign z[7:0] = inputVector[1:0];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
