
assign out = !((in1 & in2) | (in3));

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
