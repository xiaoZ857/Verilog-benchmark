
// TopModule.v
// 10‑state decade counter (1‑10 inclusive)
// Synchronous active‑high reset

module TopModule (
    input  wire        clk,    // Clock
    input  wire        reset,  // Synchronous active‑high reset
    output reg  [3:0]  q       // 4‑bit counter output
);

    // Synchronous logic
    always @(posedge clk) begin
        if (reset) begin
            q <= 4'd1;          // Reset counter to 1
        end
        else if (q == 4'd10) begin
            q <= 4'd1;          // Wrap from 10 back to 1
        end
        else begin
            q <= q + 4'd1;      // Increment counter
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
