
// TopModule.v
// 3‑bit to 16‑bit combinational lookup table
module TopModule (
    input  wire [2:0] a,          // 3‑bit address
    output reg  [15:0] q          // 16‑bit data output
);

    // Combinational logic – no clock
    always @(*) begin
        case (a)
            3'd0: q = 16'h1232;
            3'd1: q = 16'haee0;
            3'd2: q = 16'h27d4;
            3'd3: q = 16'h5a0e;
            3'd4: q = 16'h2066;
            3'd5: q = 16'h64ce;
            3'd6: q = 16'hc526;
            3'd7: q = 16'h2f19;
            default: q = 16'h0000;   // optional – covers X/unknown
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
