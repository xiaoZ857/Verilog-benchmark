

module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] pedge
);

always @(posedge clk) begin
  pedge = in;
end

always @(posedge clk) begin
  for (int i = 0; i < 8; i++) begin
    if (in[i] != pedge[i]) begin
      pedge[i] = in[i];
    end
  end
end

always @(posedge clk) begin
  for (int i = 0; i < 8; i++) begin
    if (in[i] == 0 && pedge[i] == 0) begin
      if (in[i] == 1) begin
        pedge[i] = 1;
      end
    end
  end
end

endmodule
