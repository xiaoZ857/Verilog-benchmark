
module TopModule (
  input clk,
  input load,
  input ena,
  input [1:0] amount,
  input [63:0] data,
  output reg [63:0] q
);

always @(posedge clk) begin
    if (load)
        q <= data;
    else if (ena) begin
        switch (amount)
            // Shift left by 1 bit
            (2'b00 : q <= {q[62], q[63]};
             // Shift left by 8 bits
             (2'b01 : q <= {q[71], q[64:0]});
             // Shift right by 1 bit
             (2'b10 : q <= {q[62], q[63:0]});
             // Shift right by 8 bits
             (2'b11 : begin
                 local: [64:0] temp;
                 for(int i = 0; i < 64; i++)
                     temp[i] = q[i+amount];
                 q <= temp;
             end)
        end
    end
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
