
module TopModule (
  input [15:0] in,
  output [7:0] out_hi,
  output [7:0] out_lo
);

  // Assign the upper byte of the input to out_hi
  assign out_hi = in

// VERILOG-EVAL: endmodule not found
