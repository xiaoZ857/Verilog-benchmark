
module TopModule (
  input a,
  input b,
  output out_assign,
  output reg out_alwaysblock
);

// Continuous assignment using an assign statement
assign out_assign = a & b;

// Combinational always block using @(*) for sensitivity
always @(*) begin
  out_alwaysblock = a & b;
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
