
module TopModule (
  input wire clk,
  input [7:0] in,
  output reg [7:0] pedge
);

always @(posedge clk) begin
  for (int i = 0; i < 8; i++) begin
    if (in[i] && ~pedge[i]) // if previous state was 0 and current state is 1
      pedge[i] <= 1;        // set output bit the cycle after a 0 to 1 transition occurs
    else if (!in[i] && pedge[i])
      pedge[i] <= 0;        // reset output bit when current state is 0 and previous state was 1
  end
end

initial begin
  pedge <= 0;                   // initialize all output bits to 0
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
