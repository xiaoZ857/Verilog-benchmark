
assign one = 1'b1; // Continuously assign logic high to the output

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
