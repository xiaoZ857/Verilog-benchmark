
module TopModule (
  input in,
  output out
);
// Assign the NOT operation to the output signal
assign out = ~in;

// VERILOG-EVAL: endmodule not found
