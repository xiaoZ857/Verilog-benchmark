
module TopModule (
  input cpu_overheated,
  output reg shut_off_computer,
  input arrived,
  input gas_tank_empty,
  output reg keep_driving
);
always @(*) begin
    if (cpu_overheated)
        shut_off_computer = 1'b0;  // Active low

    else 
        if (~arrived && gas_tank_empty) // If arrived and gas tank empty, don't keep driving
            keep_driving = 1'b0;
        else 
            if (arrived && ~gas_tank_empty)
                keep_driving = 1'b1;  // Keep driving as long as arrived but not empty
            else 
                shut_off_computer = 1'b1;  // Shut off computer by default
end

// VERILOG-EVAL: endmodule not found
