
module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);

  // Internal register to hold next state
  reg [255:0] next_q;
  
  integer i, j, k;
  reg [3:0] neighbor_count;
  reg current_cell;
  reg [3:0] row_above, row_below, col_left, col_right;
  reg [4:0] neighbor_idx;
  
  always @(*) begin
    // Default: keep current state
    next_q = q;
    
    // Calculate next state for each cell
    for (i = 0; i < 16; i = i + 1) begin
      for (j = 0; j < 16; j = j + 1) begin
        // Calculate wrap-around indices
        row_above = (i == 0) ? 15 : i - 1;
        row_below = (i == 15) ? 0 : i + 1;
        col_left = (j == 0) ? 15 : j - 1;
        col_right = (j == 15) ? 0 : j + 1;
        
        // Count neighbours
        neighbor_count = 0;
        
        // Top row neighbours
        neighbor_idx = row_above * 16 + col_left;
        neighbor_count = neighbor_count + q[neighbor_idx];
        neighbor_idx = row_above * 16 + j;
        neighbor_count = neighbor_count + q[neighbor_idx];
        neighbor_idx = row_above * 16 + col_right;
        neighbor_count = neighbor_count + q[neighbor_idx];
        
        // Same row neighbours (left and right)
        neighbor_idx = i * 16 + col_left;
        neighbor_count = neighbor_count + q[neighbor_idx];
        neighbor_idx = i * 16 + col_right;
        neighbor_count = neighbor_count + q[neighbor_idx];
        
        // Bottom row neighbours
        neighbor_idx = row_below * 16 + col_left;
        neighbor_count = neighbor_count + q[neighbor_idx];
        neighbor_idx = row_below * 16 + j;
        neighbor_count = neighbor_count + q[neighbor_idx];
        neighbor_idx = row_below * 16

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
