
// Define timescale outside the module
`timescale 1ns / 1ps

module TopModule (
  input clk,
  input resetn,
  input [1:0] byteena,
  input [15:0] d,
  output reg [15:0] q
);

always_ff @ (posedge clk) begin
  if (!resetn) begin
    q <= 0;
  end else begin
    // Only update the selected bytes based on byteena
    if (byteena[0]) begin
      q[7:0] <= d[7:0];
    end
    if (byteena[1]) begin
      q[15:8] <= d[15:8];
    end
  end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
