
       ab
   cd  00  01  11  10
   00 | 0 | 1 | 0 | 1 |
   01 | 1 | 0 | 1 | 0 |
   11 | 0 | 1 | 0 | 1 |
   10 | 1 | 0 | 1 | 0 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
