
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);

always @(posedge clk) begin
    if (reset) begin
        current_state <= IDLE;
        done <= 1'b0;
    end else begin
        case (current_state)
            IDLE: begin
                done <= 1'b0;
                if (in[3] == 1'b1) begin
                    current_state <= BYTE1;
                end else begin
                    current_state <= IDLE;
                end
            end
            
            BYTE1: begin
                if (in[3] == 1'b1) begin
                    // This could be byte 1 of a new message
                    current_state <= BYTE1;
                end else begin
                    current_state <= BYTE2;
                end
            end
            
            BYTE2: begin
                if (in[3] == 1'b1) begin
                    // This could be byte 1 of a new message
                    current_state <= BYTE1;
                end else begin
                    // This is byte 3, signal done
                    current_state <= BYTE3;
                end
            end
            
            BYTE3: begin
                // Signal done for one cycle
                done <= 1'b1;
                if (in[3] == 1'b1) begin
                    // This is byte 1 of next message
                    current_state <= BYTE1;
                end else begin
                    current_state <= IDLE;
                end
            end
            
            default: begin
                current_state <= IDLE;
                done <= 1'b0;
            end
        endcase
    end
end

endmodule
