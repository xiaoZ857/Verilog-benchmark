
module TopModule (
  input in,
  output out
);
assign out = in;

endmodule
