
`timescale 1ns / 1ps

module TopModule (
  input clk,
  input load,
  input [9:0] data,
  output tc
) 
{
  reg [9:0] counter;

  always @(posedge clk) begin
    if (load) begin
      counter <= data;
    end else begin
      if (counter > 0) begin
        counter <= counter - 1;
      end
    end
  end

  assign tc = (counter == 0);
}
endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
