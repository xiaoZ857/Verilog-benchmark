
assign q = ~(a ^ c) | (d ^ c);

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
