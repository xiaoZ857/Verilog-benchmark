
module TopModule (
  output one
);
 ```verilog
assign one = 1'b1;
endmodule

// VERILOG-EVAL: abnormal backticks count
