

module TopModule (
  input clk,
  input load,
  input [511:0] data,
  output reg [511:0] q
);

always @(posedge clk) begin
  if (load) begin
    q <= data;
  end else begin
    for (int i = 0; i < 512; i++) begin
      if (i == 0) begin
        q[i] <= data[i] ^ 0 ^ data[i+1];
      end else if (i == 511) begin
        q[i] <= data[i] ^ data[i-1] ^ 0;
      end else begin
        q[i] <= data[i-1] ^ data[i] ^ data[i+1];
      end
    end
  end
endmodule
