
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);
reg carry;

always @(posedge clk or posedge areset) begin
    if (areset)
        carry <=

// VERILOG-EVAL: endmodule not found
