
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);

always @(posedge clk) begin
    if (reset) begin
        current_state <= 2'b00;
    end else begin
        current_state <= next_state;
    end
end

always @(*) begin
    case (current_state)
        2'b00: begin
            if (in) next_state = 2'b01;
            else next_state = 2'b00;
        end
        2'b01: begin
            if (in) next_state = 2'b01;
            else next_state = 2'b10;
        end
        2'b10: begin
            if (in) next_state = 2'b11;
            else next_state = 2'b00;
        end
        2'b11: begin
            if (in) next_state = 2'b01;
            else next_state = 2'b10;
        end
        default: next_state = 2'b00;
    endcase
end

assign out = (current_state == 2'b11);

endmodule
