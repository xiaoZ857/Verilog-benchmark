

module TopModule (
  input [254:0] in,
  output reg [7:0] out
);



// VERILOG-EVAL: endmodule not found
