
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);
always @(*) begin
    case (y)
        3'b000, // State A
        3'b001, // State B
        3'b011, // State D
        3'b101: Y2 = w; // Transition to states C, E, F

        3'b010, // State C
        3'b100, // State E
        3'b110: Y2 = ~w; // Transition to states D, D, F

        default: Y2 = y[2]; // Remain in state F or undefined state
    endcase
end
endmodule
