
module TopModule (
    input clk,
    input reset,
    input x,
    output reg z
);

    // State register
    reg [2:0] y;
    reg [2:0] next_y;

    // Synchronous reset and state transition logic
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            y <= 3'b000; // Reset to initial state S0
            z <= 0;      // Ensure output is also reset
        end else begin
            y <= next_y;
        end
    end

    // Next state and output logic
    always @(*) begin
        case (y)
            3'b000: begin
                next_y = (x == 0) ? 3'b000 : 3'b001; // S0 -> S0 if x=0, else S1
                z = 0;
            end
            3'b001: begin
                next_y = (x == 0) ? 3'b001 : 3'b100; // S1 -> S1 if x=0, else S4
                z = 0;
            end
            3'b010: begin
                next_y = (x == 0) ? 3'b010 : 3'b001; // S2 -> S2 if x=0, else S1
                z = 0;
            end
            3'b011: begin
                next_y = (x == 0) ? 3'b001 : 3'b010; // S3 -> S1 if x=0, else S2
                z = 1;
            end
            3'b100: begin
                next_y = (x == 0) ? 3'b011 : 3'b100; // S4 -> S3 if x=0, else S4
                z = 1;
            end
            default: begin
                next_y = 3'b000; // Default case to handle unexpected states
                z = 0;
            end
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
