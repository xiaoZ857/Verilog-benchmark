
module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);
always @(posedge clk) begin
  if (reset && q == 1'b0) begin
    count <= 1;
    q <= 1'b0;
  end else begin
    // Increment the count and wrap around when it reaches 10
    count <= count + 1;
    q <= count[3:0];
  end
end

// VERILOG-EVAL: endmodule not found
