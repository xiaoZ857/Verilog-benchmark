
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);

// State encoding
parameter S0 = 1'b0;
parameter S1 = 1'b1;

reg state, next_state;

// State register with asynchronous reset
always @(posedge clk or posedge areset) begin
    if (areset)
        state <= S0;
    else
        state <= next_state;
end

// Next state logic
always @(*) begin
    case (state)
        S0: begin
            if (x)
                next_state = S1;
            else
                next_state = S0;
        end
        S1: begin
            next_state = S1;
        end
        default: next_state = S0;
    endcase
end

// Output logic (Moore machine)
assign z = (state == S0) ? x : ~x;

endmodule
