
module TopModule (
  output out
);
  out = 1'b0;
endmodule
