
module TopModule (
  input clk,
  input x,
  input [2:0] y,
  output reg Y0,
  output reg z
);


// VERILOG-EVAL: endmodule not found
