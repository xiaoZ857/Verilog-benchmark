
module TopModule (
  input a,
  input b,
  input c,
  input d,
  input e,
  output [24:0] out
);
assign out[24] = ~(a & ~b);
assign out[23] = ~(a & ~c);
assign out[22] = ~(a & ~d);
assign out[21] = ~(a & ~e);

assign out[20] = ~(b & ~a);
assign out[19] = ~(b & ~c);
assign out[18] = ~(b & ~d);
assign out[17] = ~(b & ~e);

assign out[16] = ~(c & ~a);
assign out[15] = ~(c & ~b);
assign out[14] = ~(c & ~d);
assign out[13] = ~(c & ~e);

assign out[12] = ~(d & ~a);
assign out[11] = ~(d & ~b);
assign out[10] = ~(d & ~c);
assign out[9] = ~(d & ~e);

assign out[8] = ~(e & ~a);
assign out[7] = ~(e & ~b);
assign out[6] = ~(e & ~c);
assign out[5] = ~(e & ~d);

assign out[4] = ~((~a ^ a) & (~b ^ b));
assign out[3] = ~((~a ^ a) & (~c ^ c));
assign out[2] = ~((~a ^ a) & (~d ^ d));
assign out[1] = ~((~a ^ a) & (~e ^ e));
assign out[0] = ~(a ^ b);

endmodule
