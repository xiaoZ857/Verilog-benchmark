
module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);
// State encoding
localparam OFF = 1'b0;
localparam ON  = 1'b1;

// State register
logic state, next_state;

// Sequential logic – synchronous reset
always_ff @(posedge clk) begin
    if (reset)
        state <= OFF;
    else
        state <= next_state;
end

// Next‑state logic
always_comb begin
    case (state)
        OFF: next_state = j ? ON : OFF;
        ON:  next_state = k ? OFF : ON;
        default: next_state = OFF; // safety
    endcase
end

// Moore output (same as state)
assign out = state;

endmodule
