
module TopModule(
    input clk,
    input resetn,
    input x,
    input y,
    output f,
    output g
);

reg [1:0] state; // State of the FSM (A, B, C)
reg [1:0] nextState; // Next state of the FSM
reg [1:0] prevState; // Previous state of the FSM

// Initialize states
initial begin
    state = 2'b00;
    nextState = 2'b00;
    prevState = 2'b00;
end

always @(posedge clk) begin
    if (!resetn) begin // Reset
        state <= 2'b00; // Reset to state A
        nextState <= 2'b00; // Next state is still A
        prevState <= 2'b00; // Previous state is still A
    end else begin // Not reset
        case(state)
            2'b00: // State A
                if (x == 1) begin // x = 1, move to B
                    nextState <= 2'b01;
                end else if (x == 0 && y == 1) begin // x = 0 and y = 1, set g = 1
                    g <= 1;
                    nextState <= 2'b10; // Move to C
                end else if (x == 0 && y == 0) begin // x = 0 and y = 0, stay in A
                    nextState <= 2'b00;
                end else begin // Invalid input, stay in A
                    nextState <= 2'b00;
                end
        endcase

        case(nextState)
            2'b01: // State B
                if (x == 1) begin // x = 1, move to C
                    nextState <= 2'b10;
                end else if (x == 0 && y == 1) begin // x = 0 and y = 1, set g = 1
                    g <= 1;
                    nextState <= 2'b11; // Move to D
                end else if (x == 0 && y == 0) begin // x = 0 and y = 0, move back to A
                    nextState <= 2'b00;
                end else begin // Invalid input, move back to B
                    nextState <= 2'b01;
                end

            2'b10: // State C
                if (x == 1) begin // x = 1, set g = 0 and move to A
                    f <= 1;
                    g <= 0;
                    nextState <= 2'b00;
                end else if (y == 1 && prevState == 2'b01) begin // y = 1 and previous state was B, set g = 1
                    g <= 1;
                    nextState <= 2'b11; // Move to D
                end else if (x == 0 && y == 0) begin // x = 0 and y = 0, move back to A
                    nextState <= 2'b00;
                end else begin // Invalid input, set g = 0 and stay in C
                    f <= 1;
                    g <= 0;
                    nextState <= 2'b10;
                end

            2'b11: // State D
                if (y == 1) begin // y = 1, move back to A
                    f <= 1;
                    g <= 0;
                    nextState <= 2'b00;
                end else if (x == 0 && prevState == 2'b10) begin // x = 0 and previous state was C, set g = 0
                    g <= 0;
                    nextState <= 2'b01; // Move back to B
                end else begin // Invalid input, move back to D
                    f <= 1;
                    g <= 0;
                    nextState <= 2'b11;
                end

        endcase

        prevState <= state; // Update previous state
    end
endmodule

// VERILOG-EVAL: errant inclusion of module definition
