
module TopModule (
    input  wire clk,    // clock
    input  wire j,      // input that drives OFF → ON transition
    input  wire k,      // input that drives ON  → OFF transition
    input  wire reset,  // active‑high synchronous reset
    output wire out     // Moore output (same as state)
);

    // State

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
