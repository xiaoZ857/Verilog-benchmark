

module TopModule (
  input [4:1] x,
  output logic f
);

always_ff @(posedge clk) begin
    case (x)
        4'b0100, 4'b0110, 4'b1000, 4'b1010, 4'b1100, 4'b1110: f <= 1;
        4'b0010, 4'b0101, 4'b1001, 4'b1011: f <= 0;
        default: f <= 1; // Use don't-care to output 1
    endcase
end

endmodule
