
module TopModule (
    input [99:0] a,
    input [99:0] b,
    input sel,
    output reg [99:0] out
);

  // Assign the output based on the select signal
  always @(*) begin
    if (sel == 1'b0)
      out = a;
    else
      out = b;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
