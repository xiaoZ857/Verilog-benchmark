
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);
always @(*) begin
    case (y)
        3'b000, // State A
        3'b001, // State B, transition on w=0 to C
        3'b011: Y2 = ~w; // States D and E transition on w=1 back to A
        
        3'b010, // State C
        3'b100: Y2 = 1'b0; // State F

        default: Y2 = 1'bx;
    endcase
end
endmodule
