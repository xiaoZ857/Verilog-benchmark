
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

// State encoding
parameter WALK_LEFT = 3'd0;
parameter WALK_RIGHT = 3'd1;
parameter FALL_LEFT = 3'd2;
parameter FALL_RIGHT = 3'd3;
parameter DIG_LEFT = 3'd4;
parameter DIG_RIGHT = 3'd5;

reg [2:0] state, next_state;

// State transition logic
always @(*) begin
    next_state = state;
    
    case (state)
        WALK_LEFT: begin
            // Fall has highest priority
            if (!ground) begin
                next_state = FALL_LEFT;
            end
            // Dig has second priority
            else if (dig) begin
                next_state = DIG_LEFT;
            end
            // Direction change has lowest priority
            else if (bump_left || bump_right) begin
                next_state = WALK_RIGHT;
            end
        end
        
        WALK_RIGHT: begin
            // Fall has highest priority
            if (!ground) begin
                next_state = FALL_RIGHT;
            end
            // Dig has second priority
            else if (dig) begin
                next_state = DIG_RIGHT;
            end
            // Direction change has lowest priority
            else if (bump_left || bump_right) begin
                next_state = WALK_LEFT;
            end
        end
        
        FALL_LEFT: begin
            if (ground) begin
                next_state = WALK_LEFT;
            end
        end
        
        FALL_RIGHT: begin
            if (ground) begin
                next_state = WALK_RIGHT;
            end
        end
        
        DIG_LEFT: begin
            if (!ground) begin
                next_state = FALL_LEFT;
            end
        end
        
        DIG_RIGHT: begin
            if (!ground) begin
                next_state = FALL_RIGHT;
            end
        end
    endcase
end

// State register
always @(posedge clk or posedge areset) begin
    if (areset) begin
        state <= WALK_LEFT;
    end else begin
        state <= next_state;
    end
end

// Output logic (Moore machine)
assign walk_left = (state == WALK_LEFT);
assign walk_right = (state == WALK_RIGHT);
assign aaah = (state == FALL_LEFT) || (state == FALL_RIGHT);
assign digging = (state == DIG_LEFT) || (state == DIG_RIGHT);

endmodule
