
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);

// FSM for serial data reception with start/stop bits
reg [2:0] state, next_state;
reg [7:0] data_reg;
reg [2:0] bit_count;
reg done_reg;

// State definitions
localparam IDLE = 3'd0;
localparam START = 3'd1;
localparam DATA = 3'd2;
localparam STOP = 3'd3;
localparam WAIT_STOP = 3'd4;

// State register
always @(posedge clk) begin
    if (reset) begin
        state <= IDLE;
        data_reg <= 8'b0;
        bit_count <= 3'b0;
        done_reg <= 1'b0;
    end else begin
        state <= next_state;
        
        case (state)
            START: begin
                data_reg <= 8'b0;
                bit_count <= 3'b0;
                done_reg <= 1'b0;
            end
            DATA: begin
                // Shift in data bits (LSB first)
                data_reg <= {data_reg[6:0], in};
                bit_count <= bit_count + 1;
                done_reg <= 1'b0;
            end
            STOP: begin
                if (in == 1) begin
                    done_reg <= 1'b1;
                end else begin
                    done_reg <= 1'b0;
                end
            end
            WAIT_STOP: begin
                if (in == 1) begin
                    done_reg <= 1'b1;
                end else begin
                    done_reg <= 1'b0;
                end
            end
            default: begin
                done_reg <= 1'b0;
            end
        endcase
    end
end

// Next state logic
always @(*) begin
    next_state = state;
    case (state)
        IDLE: begin
            if (in == 0) begin
                next_state = START;
            end
        end
        START: begin
            next_state = DATA;
        end
        DATA: begin
            if (bit_count == 3'd7) begin
                next_state = STOP;
            end
        end
        STOP: begin
            if (in == 1) begin
                next_state = IDLE;
            end else begin
                next_state = WAIT_STOP;
            end
        end
        WAIT_STOP: begin
            if (in == 1) begin
                next_state = IDLE;
            end
        end
    endcase
end

// Output assignments
assign out_byte = data_reg;
assign done = done_reg;

endmodule
