
module TopModule (
  input clk,
  input d,
  input ar,
  output logic q
);
always @(posedge clk) begin
  if (ar)
    q <= 1'b0;
  else
    q <= d;
endmodule
