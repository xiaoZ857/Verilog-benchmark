
//=====================================================================
//  TopModule
//  Recognises 8‑bit keyboard scancodes for the keys 0–9.
//  If the input matches one of the 10 codes, it outputs the key value
//  (0‑9) on `out` and sets `valid` to 1.  Otherwise both outputs are 0.
//=====================================================================
module TopModule (
    input  wire [7:0] code,   // 8‑bit scancode from the keyboard
    output reg  [3:0] out,    // 4‑bit key value (0‑9)
    output reg        valid   // 1 if a valid key was detected
);

    // Combinational logic – no clock needed
    always @(*) begin
        // Default: no key recognised
        out   = 4'd0;
        valid = 1'b0;

        // Map each recognised scancode to its key value
        case (code)
            8'h45: begin out = 4'd0; valid = 1'b1; end
            8'h16: begin out = 4'd1; valid = 1'b1; end
            8'h1e: begin out = 4'd2; valid = 1'b1; end
            8'h26: begin out = 4'd3; valid = 1'b1; end
            8'h25: begin out = 4'd4; valid = 1'b1; end
            8'h2e: begin out = 4'd5; valid = 1'b1; end
            8'h36: begin out = 4'd6; valid = 1'b1; end
            8'h3d: begin out = 4'd7; valid = 1'b1; end
            8'h3e: begin out = 4'd8; valid = 1'b1; end
            8'h46: begin out = 4'd9; valid = 1'b1; end
            default: ; // already set to 0/0
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
