
module TopModule (
  input [6:1] y,
  input w,
  output Y2,
  output Y4
);
always @(posedge clk) begin
  if (y[6] || y[5]) Y2 <= 0'b0;            // A or B -> Y2 = 0
  else if (y[3]) Y2 <= 1'b1;               // C -> Y2 = 1
  else if (y[4]) Y2 <= y[6];              // D -> Y2 = A
  else if (y[2]) Y2 <= y[0];              // E -> Y2 = A
  else if (y[1]) Y2 <= y[3];              // F -> Y2 = C
end

always @(posedge clk) begin
  if (y[6]) Y4 <= 0'b0;                // A -> Y4 = 0
  else if (y[5]) Y4 <= y[4];           // B -> Y4 = D
  else if (y[3]) Y4 <= y[2];           // C -> Y4 = E
  else if (y[4]) Y4 <= w;              // D -> Y4 = w
  else if (y[2]) Y4 <= y[5];           // E -> Y4 = B
  else if (y[1]) Y4 <= y[6];           // F -> Y4 = A
end

// Add `timescale` directive outside the module definition
`timescale 1ns / 1ps

// VERILOG-EVAL: endmodule not found
