
module TopModule (
    input [99:0] in,
    output reg [99:0] out
);

always @(posedge clk)
begin
    for (int i = 0; i < 100; i++)
        out[i] <= in[99-i];
end

// Assuming a clock signal 'clk' is provided externally.
// If not provided, replace "@(posedge clk)" with "@" to make it edge-triggered on positive or negative transition.

endmodule

// VERILOG-EVAL: errant inclusion of module definition
