
module TopModule (
  input a,
  input b,
  output out
);
// Define the XNOR gate module
module XNORGate(
    // Inputs
    input a, 
    input b, 
    // Output
    output out
);

    // Assign the output based on the inputs
    assign out = !((a & b) | (~a & ~b));

endmodule

// Define the TopModule that includes the XNOR gate
module TopModule(
    // Inputs
    input a, 
    input b,
    // Output
    output out
);

    // Instantiate the XNOR gate module
    XNORGate xnor_gate (
        .a(a),
        .b(b),
        .out(out)
    );

endmodule

// VERILOG-EVAL: errant inclusion of module definition
