
module TopModule (
  input [2:0] vec,
  output [2:0] outv,
  output o2,
  output o1,
  output o0
);
Here's the implementation of the `TopModule` in Verilog, as per the given description:

---

### ✅ **Module Overview**

- **Inputs**: A 3-bit vector `vec`.
- **Outputs**:
  - A 3-bit

// VERILOG-EVAL: endmodule not found
