
module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);

  wire carry0, carry1, carry2, carry3;
  
  // First full adder (LSB)
  assign sum[0] = x[0] ^ y[0] ^ 1'b0;
  assign carry0 = (x[0] & y[0]) | (x[0] & 1'b0) | (y[0] & 1'b0);
  
  // Second full adder
  assign sum[1] = x[1] ^ y[1] ^ carry0;
  assign carry1 = (x[1] & y[1]) | (x[1] & carry0) | (y[1] & carry0);
  
  // Third full adder
  assign sum[2] = x[2] ^ y[2] ^ carry1;
  assign carry2 = (x[2] & y[2]) | (x[2] & carry1) | (y[2] & carry1);
  
  // Fourth full adder (MSB)
  assign sum[3] = x[3] ^ y[3] ^ carry2;
  assign carry3 = (x[3] & y[3]) | (x[3] & carry2) | (y[3] & carry2);
  
  // Overflow bit (final carry out)
  assign sum[4] = carry3;
  
endmodule
