
module TopModule (
  input [7:0] in,
  output reg [2:0] pos
);

always @(*) begin
  if (in[0]) begin
    pos = 3'b000;
  end else if (in[1]) begin
    pos = 3'b001;
  end else if (in[2]) begin
    pos = 3'b010;
  end else if (in[3]) begin
    pos = 3'b011;
  end else if (in[4]) begin
    pos = 3'b100;
  end else if (in[5]) begin
    pos = 3'b101;
  end else if (in[6]) begin
    pos = 3'b110;
  end else if (in[7]) begin
    pos = 3'b111;
  end else begin
    pos = 3'b000; // Default to zero if no bits are high
  end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
