
typedef enum State { A, B, C, D } State;

module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
    State current_state = A;
    
    always @(posedge clk) begin
        if (reset) begin
            current_state <= A;
        end else begin
            case (current_state)
                A: 
                    case (in)
                        0: current_state <= A;
                        1: current_state <= B;
                    endcase
                B:
                    case (in)
                        0: current_state <= C;
                        1: current_state <= B;
                    endcase
                C:
                    case (in)
                        0: current_state <= A;
                        1: current_state <= D;
                    endcase
                D:
                    case (in)
                        0: current_state <= C;
                        1: current_state <= B;
                    endcase
            endcase
        end
    end
    
    always @(*) begin
        case (current_state)
            A: out = 0;
            B: out = 0;
            C: out = 0;
            D: out = 1;
        endcase
    end
endmodule

// VERILOG-EVAL: errant inclusion of module definition
