
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
// State transition logic
always @(*) begin
    case (current_state)
        A: next_state = (w == 0) ? B : A;
        B: next_state = (w == 0) ? C : D;
        C: next_state = (w == 0) ? E : D;
        D: next_state = (w == 0) ? F : A;
        E: next_state = (w == 1) ? D : E; // Corrected condition
        F: next_state = (w == 0) ? C : D; // Corrected condition
        default: next_state = A;
    endcase
end

// Output logic
always @(*) begin
    case (current_state)
        E: z = w; // Output based on state E and input w
        F: z = ~w; // Output based on state F and inverted input w
        default: z = 0;  // Default output value
    endcase
end

// State update logic remains unchanged
always @(posedge clk or posedge reset) begin
    if (reset)
        current_state <= A;
    else
        current_state <= next_state;
end

endmodule
