
module TopModule (
  input a,
  input b,
  output out
);
assign out = a ^ b; endmodule

// VERILOG-EVAL: endmodule not found
