
module TopModule (
  input in,
  input [1:0] state,
  output reg [1:0] next_state,
  output out
);
// Output logic – Moore output depends only on the current state
assign out = (state == 2'b11);   // 1 only in state D, 0 otherwise

// Combinational logic for next state
always_comb begin
  case (state)
    2'b00: begin // State A
      next_state = (in == 1'b0) ? 2'b00 : 2'b01; // stay A or go to B
    end
    2'b01: begin // State B
      next_state = (in == 1'b0) ? 2'b10 : 2'b01; // go to C or stay B
    end
    2'b10: begin // State C
      next_state = (in == 1'b0) ? 2'b00 : 2'b11; // go to A or D
    end
    2'b11: begin // State D
      next_state = (in == 1'b0) ? 2'b10 : 2'b01; // go to C or B
    end
    default: begin
      next_state = 2'b00; // safe default
    end
  endcase
end

endmodule
