
module TopModule (
  input mode,
  input too_cold,
  input too_hot,
  input fan_on,
  output heater,
  output aircon,
  output fan
);

  // Heater control logic
  assign heater = mode & too_cold;
  
  // Air conditioner control logic
  assign aircon = ~mode & too_hot;
  
  // Fan control logic - turns on when heater or AC is on, or when user requests it
  assign fan = heater | aircon | fan_on;

endmodule
