

module TopModule (
  input [1023:0] in,
  input [7:0] sel,
  output [3:0] out
);

reg [3:0] out_reg;

always @(posedge clk) begin
    case (sel)
        8'b00000000: out_reg <= in[3:0];
        8'b00000001: out_reg <= in[7:4];
        8'b00000010: out_reg <= in[11:8];
        8'b00000011: out_reg <= in[15:12];
        8'b00000100: out_reg <= in[19:16];
        8'b00000101: out_reg <= in[23:20];
        8'b00000110: out_reg <= in[27:24];
        8'b00000111: out_reg <= in[31:28];
        8'b00001000: out_reg <= in[35:32];
        8'b00001001: out_reg <= in[39:36];
        8'b00001010: out_reg <= in[43:40];
        8'b00001011: out_reg <= in[47:44];
        8'b00001100: out_reg <= in[51:48];
        8'b00001101: out_reg <= in[55:52];
        8'b00001110: out_reg <= in[59:56];
        8'b00001111: out_reg <= in[63:60];
        8'b00010000: out_reg <= in[67:64];
        8'b00010001: out_reg <= in[71:68];
        8'b00010010: out_reg <= in[75:72];
        8'b00010011: out_reg <= in[79:76];
        8'b00010100: out_reg <= in[83:80];
        8'b00010101: out_reg <= in[87:84];
        8'b00010110: out_reg <= in[91:88];
        8'b00010111: out_reg <= in[95:92];
        8'b00011000: out_reg <= in[99:96];
        8'b00011001: out_reg <= in[103:100];
        8'b00011010: out_reg <= in[107:104];
        8'b00011011: out_reg <= in[111:108];
        8'b00011100: out_reg <= in[115:112];
        8'b00011101: out_reg <= in[119:116];
        8'b00011110: out_reg <= in[123:120];
        8'b00011111: out_reg <= in[127:124];
        8'b00100000: out_reg <= in[131:128];
        8'b00100001: out_reg <= in[135:132];
        8'b00100010: out_reg <= in[139:136];
        8'b00100011: out_reg <= in[143:140];
        8'b00100100: out_reg <= in[147:144];
        8'b00100101: out_reg <= in[151:148];
        8'b00100110: out_reg <= in[155:152];
        8'b00100111: out_reg <= in[159:156];
        8'b00101000: out_reg <= in[163:160];
        8'b00101001: out_reg <= in[167:164];
        8'b00101010: out_reg <= in[171:168];
        8'b00101011: out_reg <= in[175:172];
        8'b00101100: out_reg <= in[179:176];
        8'b00101101: out_reg <= in[183:180];
        8'b00101110: out_reg <= in[187:184];
        8'b00101111: out_reg <= in[191:188];
        8'b00110000: out_reg <= in[195:192];
        8'b00110001: out_reg <= in[199:196];
        8'b00110010: out_reg <= in[203:200];
        8'b00110011: out_reg <= in[207:204];
        8'b00110100: out_reg <= in[211:208];
        8'b00110101: out_reg <= in[215:212];
        8'b00110110: out_reg <= in[219:216];
        8'b00110111: out_reg <= in[223:220];
        8'b00111000: out_reg <= in[227:224];
        8'b00111001: out_reg <= in[231:228];
        8'b00111010: out_reg <= in

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
