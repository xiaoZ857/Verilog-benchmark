
assign out_hi = in[15:8];
assign out_lo = in[7:0];

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
