
module TopModule (
  input [7:0] in,
  output parity
);
always @(posedge clk) begin
  if (clk == 1'b0) // Reset condition
    parity <= 1'b1; // Initialize parity as '1'
  else // Normal operation
    parity ^= in; // XOR all input bits with the current parity value
end

always @(negedge clk) begin
  if (clk == 1'b0) // Reset condition
    $display("Parity: %b", parity); // Dump initial parity value
end

initial begin
  $dumpfile("parity_checker.vcd");
  $dumpvars(0, TopModule);
  #100; // Simulation time for 100 ns
  clk = 1'b0; // Reset clock to low state
  #50; // Delay for 50 ns
  clk = 1'b1; // Set clock to high state
  repeat(8) begin
    #25; // Delay for 25 ns between each input change
    in <= in + 1; // Increment the input byte by 1 every 25 ns
  end
  #100; // Simulation time for 100 ns after the last input change
end

// VERILOG-EVAL: endmodule not found
