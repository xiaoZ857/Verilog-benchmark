
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);
  reg [2:0] state, next_state;
  
  // State encoding
  localparam S0 = 3'b000,
             S1 = 3'b001,
             S2 = 3'b010,
             S3 = 3'b011,
             S4 = 3'b100;
  
  // State register
  always @(posedge clk) begin
    if (reset)
      state <= S0;
    else
      state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      S0: next_state = data ? S1 : S0;
      S1: next_state = data ? S2 : S0;
      S2: next_state = data ? S2 : S3;
      S3: next_state = data ? S4 : S0;
      S4: next_state = S4; // stay until reset
      default: next_state = S0;
    endcase
  end
  
  // Output logic
  assign start_shifting = (state == S4);

endmodule
