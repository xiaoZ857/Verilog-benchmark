
module TopModule (
  input wire clk,
  input wire j,
  input wire k,
  input wire areset,
  output reg out
);

  // State encoding
  typedef enum logic [1:0] {
    OFF = 2'b00,
    ON  = 2'b01
  } state_t;

  // Declare state register
  state_t current_state, next_state;

  // Output logic based on the current state (Moore machine)
  always @(*) begin
    case(current_state)
      OFF: out = 0;
      ON : out = 1;
      default: out = 0; // Default case for safety
    endcase
  end

  // Next state logic and synchronous reset handling
  always_ff @(posedge clk or posedge areset) begin
    if (areset) begin
      current_state <= OFF; // Asynchronous reset to OFF
    end else begin
      current_state <= next_state;
    end
  end

  // Next state logic based on the current state and inputs j, k
  always @(*) begin
    case(current_state)
      OFF: begin
        if (j) 
          next_state = ON;
        else 
          next_state = OFF;
      end
      
      ON : begin
        if (k) 
          next_state = OFF;
        else 
          next_state = ON;
      end
      
      default: next_state = OFF; // Default case for safety
    endcase
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
