
module TopModule (
  input [7:0] code,
  output reg [3:0] out,
  output reg valid
);
assign out = $signed(code[6:1]) == 8'h45 ? 4'd0 : 
               $signed(code[6:1]) == 8'h16 ? 4'd1 : 
               $signed(code[6:1]) == 8'h1e ? 4'd2 : 
               $signed(code[6:1]) == 8'h26 ? 4'd3 : 
               $signed(code[6:1]) == 8'h25 ? 4'd4 : 
               $signed(code[6:1]) == 8'h2e ? 4'd5 : 
               $signed(code[6:1]) == 8'h36 ? 4'd6 : 
               $signed(code[6:1]) == 8'h3d ? 4'd7 : 
               $signed(code[6:1]) == 8'h3e ? 4'd8 : 
               $signed(code[6:1]) == 8'h46 ? 4'd9 : 
               4'd0, valid = 1'b0;

always @(posedge clk) begin
    if (code[7] == 1'b1 && code[6] == 1'b0 && code[5] == 1'b0 && code[4] == 1'b0 && code[3] == 1'b0 && code[2] == 1'b0 && code[1] == 1'b0 && code[0] == 1'b0)
        valid = 1'b1;
    else
        valid = 1'b0;
end

// VERILOG-EVAL: endmodule not found
