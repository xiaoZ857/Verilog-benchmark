
// 7458 – 4 AND gates + 2 OR gates
// p1y  = (p1a & p1b & p1c) | (p1d & p1e & p1f)
// p2y  = (p2a & p2b)       | (p2c & p2d)

module TopModule (
    input  p1a, p1b, p1c, p1d, p1e, p1f,   // 6 inputs for the first OR
    output p1y,                              // 1st OR output
    input  p2a, p2b, p2c, p2d,              // 4 inputs for the second OR
    output p2y                               // 2nd OR output
);

    // 3‑input ANDs for the first OR
    wire and1 = p1a & p1b & p1c;
    wire and2 = p1d & p1e & p1f;

    // 2‑input ANDs for the second OR
    wire and3 = p2a & p2b;
    wire and4 = p2c & p2d;

    // OR the results
    assign p1y = and1 | and2;
    assign p2y = and3 | and4;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
