
module TopModule (
  input clk,
  input resetn,
  input [1:0] byteena,
  input [15:0] d,
  output reg [15:0] q
);
  reg [15:0] dff_q [0:15];

  always @(posedge clk or negedge resetn) begin
    if (!resetn) begin
      q <= 0;
      for (integer i = 0; i < 16; i = i + 1) begin
        dff_q[i] <= 0;
      end
    end else begin
      // Update the flip-flops based on byteena
      if (byteena[1]) begin
        q[15:8] <= d[15:8];
      end
      if (byteena[0]) begin
        q[7:0] <= d[7:0];
      end
    end
  end
endmodule
