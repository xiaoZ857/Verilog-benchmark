
module TopModule (
  input clk,
  input reset,
  input ena,
  output reg pm,
  output reg [7:0] hh,
  output reg [7:0] mm,
  output reg [7:0] ss
);
always @(posedge clk or posedge reset) begin
    if (reset) begin
        {pm, hh, mm, ss} <= 12'b000000010110; // Reset to "12:00 AM"
    end else if (ena) begin
        // Update seconds
        if (ss == 8'd59) begin
            ss <= 8'd0;
            // Update minutes
            if (mm == 8'd59) begin
                mm <= 8'd0;
                // Update hours and pm
                if (hh == 8'd12) begin
                    hh <= 8'd1;
                    pm <= ~pm;
                end else if (hh == 8'd11) begin
                    hh <= 8'd12;
                end else begin
                    hh <= hh + 1;
                end
            end else begin
                mm <= mm + 1;
            end
        end else begin
            ss <= ss + 1;
        end
    end
end
endmodule
