
module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);
reg state;

always @(posedge clk or negedge aresetn) begin
  if (!aresetn) begin
    state <= 0;
    z <= 0;
  end else begin
    case (state)
      0: begin
        if (x == 1)
          state <= 1;
        else
          state <= 0;
        z <= 0;
      end
      1: begin
        if (x == 0)
          state <= 2;
        else
          state <= 1;
        z <= 0;
      end
      2: begin
        if (x == 1)
          state <= 1;
        else
          state <= 0;
        z <= 1;
      end
    endcase
  end
endmodule
