
module TopModule(
    input a, // Present for 55ns to 90ns period
    input b,
    input c,
    input d,
    output q
);

    always @(*)
        q <= (c & ~d) | (~a & ~b);
endmodule

// VERILOG-EVAL: errant inclusion of module definition
