
module TopModule (
  input clk,
  input reset,
  output [3:1] ena,
  output reg [15:0] q
);


// VERILOG-EVAL: endmodule not found
