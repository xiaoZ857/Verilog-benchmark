
module TopModule (
  input clk,
  input reset,
  input x,
  output reg z
);
assign z = (reset) ? 1'b0 : ($signed<2{(x+1)/2}}[3:0]==$signed{y[1:y]}[2:y]) ^ $signed<2{((x+1)/2}>>[1]}[2:y];
always @(posedge clk or reset) begin
    if (reset)
        y <= 3'b000;
    else
        case(y)
            3'b000 : y <= 3'b001;      // y[1:0] = 00, y[2] = 0
            3'b001 : y <= 3'b010;      // y[1:0] = 01, y[2] = 0
            3'b010 : y <= 3'b001;      // y[1:0] = 10, y[2] = 0
            3'b011 : y <= 3'b000;      // y[1:0] = 11, y[2] = 0
            3'b100 : y <= 3'b110;      // y[1:0] = 01, y[2] = 1
            3'b101 : y <= 3'b001;      // y[1:0] = 10, y[2] = 1
            default:                  // y[1:0] = 00, y[2] = 1
                y <= 3'b010;
        endcase

        z <= $signed<2{(x+1)/2}}[4:y];
endmodule
