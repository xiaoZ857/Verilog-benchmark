
module TopModule (
  input d,
  input done_counting,
  input ack,
  input [9:0] state, // 10-bit one-hot current state
  output B3_next,
  output S_next,
  output S1_next,
  output Count_next,
  output Wait_next,
  output done,
  output counting,
  output shift_ena
);
assign S_next = (state[0] & ~d) | (state[1] & ~d) | (state[3] & ~d) | (state[9] & ack);
assign S1_next = (state[0] & d) | (state[1] & d);
assign B3_next = state[6];
assign Count_next = (state[7] & ~done_counting) | (state[7] & done_counting);
assign Wait_next = (state[7] & done_counting) | (state[8] & ~ack);

assign shift_ena = state[4] | state[5] | state[6] | state[7];
assign counting = state[7];
assign done = state[8];

endmodule
