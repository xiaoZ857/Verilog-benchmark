
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
// Define states using parameters
parameter A = 2'b00, B = 2'b01, C = 2'b10, D = 2'b11;

reg [1:0] current_state, next_state;

// State transition logic (combinational)
always @(*) begin
    case (current_state)
        A: next_state = in ? B : A;
        B: next_state = in ? B : C;
        C: next_state = in ? D : A;
        D: next_state = in ? B : C;
        default: next_state = A;
    endcase
end

// State register with asynchronous reset
always @(posedge clk, posedge areset) begin
    if (areset) current_state <= A;
    else current_state <= next_state;
end

// Output logic (Moore: output depends only on current state)
assign out = (current_state == D) ? 1'b1 : 1'b0;

endmodule
