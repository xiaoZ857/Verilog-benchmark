

module TopModule (
  input clk,
  input areset,
  input x,
  output z
);

  reg [1:0] state;
  reg z_reg;

  always @(posedge clk or posedge areset) begin
    if (areset) begin
      state <= 2'b00; // State A
      z_reg <= 0;
    end else begin
      case (state)
        2'b00: begin // State A
          if (x) begin
            state <= 2'b01; // Go to state B
            z_reg <= 1;
          end else begin
            state <= 2'b00; // Stay in state A
            z_reg <= 0;
          end
        end
        2'b01: begin // State B
          if (x) begin
            state <= 2'b01; // Stay in state B
            z_reg <= 0;
          end else begin
            state <= 2'b01; // Stay in state B
            z_reg <= 1;
          end
        end
        default: begin
          state <= 2'b00;
          z_reg <= 0;
        end
      endcase
    end
  end

  assign z = z_reg;

endmodule
