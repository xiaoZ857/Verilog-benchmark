
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);
always_comb begin : statesLogic
  // Walking direction
  if (cur_state == IDLE || cur_state == WALKING_LEFT) {
    walk_left <= 1; walk_right <= 0;
  } else if (cur_state == WALKING_RIGHT) {
    walk_left <= 0; walk_right <= 1;
  } else if (cur_state == FALLING || cur_state == OBSTACLE_LEFT) {
    walk_left <= 0; walk_right <= 1;
  } else if (cur_state == DIGGING_LEFT || cur_state == WALKING_RIGHT) {
    walk_left <= 1; walk_right <= 0;
  } else if (cur_state == DIGGING_RIGHT || cur_state == OBSTACLE_RIGHT) {
    walk_left <= 1; walk_right <= 0;
  } else {
    // No change in walking direction
    walk_left <= (cur_state != OBSTACLE_LEFT)? 0: walk_left;
    walk_right <= (cur_state != OBSTACLE_RIGHT)? 1: walk_right;
  }

  // AAah!
  if ((ground == 0 && dig == 0) || (bump_left && !dig && cur_state != OBSTACLE_LEFT) ||
      (bump_right && !dig && cur_state != OBSTACLE_RIGHT)) {
    aaah <= 1; digging <= 0;
  } else {
    aaah <= 0; digging <= 1;
  }

  // Digging
  if (cur_state == DIGGING_LEFT || cur_state == DIGGING_RIGHT) {
    digging <= 1;
  }
end

// Moore state machine
always @(posedge clk or negedge areset) begin : updateState
  if (areset) {
    cur_state = IDLE;
  } else {
    states_t next_state = getNextState(cur_state, bump_left, bump_right, ground, dig);
    if (next_state != cur_state) {
      cur_state = next_state;
    }
  }
end

// VERILOG-EVAL: endmodule not found
