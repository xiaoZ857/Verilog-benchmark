
module TopModule (
  input [7:0] a,
  input [7:0] b,
  output [7:0] s,
  output overflow
);
always @(posedge clk) begin
    // 2's complement addition with carry propagation and borrow generation
    s[0] <= a[0] ^ b[0] ^ carry_in;
    s[7:1] <= {a[7:1], b[7:1]} + {carry_in, carry_out} + (s[0] << 8);

    // Initialize carry-in to zero for the first addition
    if(initial_state) begin
        carry_in <= 0;
    end

    // Carry out of the MSB is carried over to next clock cycle as it's not immediately available
    assign carry_out = s[7];

    // Check for overflow based on the MSB and carry-out from the addition
    assign overflow = ~a[7] & ~b[7] | a[7] & b[7] | (carry_out && ~s[7]);
end
endmodule
