
module TopModule (
  input clk,
  input load,
  input [511:0] data,
  output reg [511:0] q
);
always @(posedge clk) begin
  if (load) begin
    q <= data;
  end else begin
    for (int i = 0; i < 512; i++) begin
      logic left = (i > 0) ? q[i-1] : 1'b0;
      logic right = (i < 511) ? q[i+1] : 1'b0;
      
      if (q[i] == 1'b1) begin
        if (left == 1'b1 && q[i] == 1'b1 && right == 1'b1)
          q[i] <= 1'b0;
        else if (left == 1'b1 && q[i] == 1'b1 && right == 1'b0)
          q[i] <= 1'b1;
        else if (left == 1'b1 && q[i] == 1'b0 && right == 1'b1)
          q[i] <= 1'b1;
        else if (left == 1'b1 && q[i] == 1'b0 && right == 1'b0)
          q[i] <= 1'b0;
        else if (left == 1'b0 && q[i] == 1'b1 && right == 1'b1)
          q[i] <= 1'b1;
        else if (left == 1'b0 && q[i] == 1'b1 && right == 1'b0)
          q[i] <= 1'b1;
        else if (left == 1'b0 && q[i] == 1'b0 && right == 1'b1)
          q[i] <= 1'b1;
        else
          q[i] <= 1'b0;
      end else begin
        if (left == 1'b1 && q[i] == 1'b1 && right == 1'b1)
          q[i] <= 1'b0;
        else if (left == 1'b1 && q[i] == 1'b1 && right == 1'b0)
          q[i] <= 1'b1;
        else if (left == 1'b1 && q[i] == 1'b0 && right == 1'b1)
          q[i] <= 1'b1;
        else if (left == 1'b1 && q[i] == 1'b0 && right == 1'b0)
          q[i] <= 1'b0;
        else if (left == 1'b0 && q[i] == 1'b1 && right == 1'b1)
          q[i] <= 1'b1;
        else if (left == 1'b0 && q[i] == 1'b1 && right == 1'b0)
          q[i] <= 1'b1;
        else if (left == 1'b0 && q[i] == 1'b0 && right == 1'b1)
          q[i] <= 1'b1;
        else
          q[i] <= 1'b0;
      end
    end
  end
endmodule
