
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);

reg [2:0] state, next_state;
reg start_shifting_reg;

parameter S0 = 3'b000;
parameter S1 = 3'b001;
parameter S2 = 3'b010;
parameter S3 = 3'b011;
parameter S4 = 3'b100;

always @(posedge clk) begin
    if (reset) begin
        state <= S0;
        start_shifting_reg <= 1'b0;
    end else begin
        state <= next_state;
        if (next_state == S4) begin
            start_shifting_reg <= 1'b1;
        end
    end
end

always @(*) begin
    case (state)
        S0: next_state = (data == 1'b1) ? S1 : S0;
        S1: next_state = (data == 1'b1) ? S2 : S0;
        S2: next_state = (data == 1'b0) ? S3 : S2;
        S3: next_state = (data == 1'b1) ? S4 : S0;
        S4: next_state = S4;
        default: next_state = S0;
    endcase
end

assign start_shifting = start_shifting_reg;

endmodule
