

module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);



// VERILOG-EVAL: endmodule not found
