
module TopModule (
  input c,
  input d,
  output [3:0] mux_in
);
 ```verilog
reg [3:0] mux_in;

always @(posedge clk or negedge a or negedge b) begin
    if (a == 0 && b == 0)
        mux_in[0] = c;
    else if (a == 1 && b == 0)
        mux_in[1] = c;
    else if (a == 1 && b == 1)
        mux_in[2] = c;
    else // a == 0 && b == 1
        mux_in[3] = c;
end

assign mux_out = {mux_in[0], mux_in[1], mux_in[2], mux_in[3]}; // 4-to-1 multiplexer output
endmodule

// VERILOG-EVAL: abnormal backticks count
