
module TopModule (
  input in1,
  input in2,
  output logic out
);


// VERILOG-EVAL: endmodule not found
