
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);
logic [2:0] state, next_state;
logic [7:0] byte1, byte2, byte3;
logic valid_byte1, valid_byte2, valid_byte3;

always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        state <= 3'b000;
        byte1 <= 8'h00;
        byte2 <= 8'h00;
        byte3 <= 8'h00;
        valid_byte1 <= 1'b0;
        valid_byte2 <= 1'b0;
        valid_byte3 <= 1'b0;
    end else begin
        state <= next_state;
        if (valid_byte1) byte1 <= in;
        if (valid_byte2) byte2 <= in;
        if (valid_byte3) byte3 <= in;
    end
end

always_comb begin
    done = 1'b0;
    out_bytes = 24'h000000;

    case (state)
        3'b000: next_state = (in[3]) ? 3'b001 : 3'b000;
        3'b001: next_state = 3'b010;
        3'b010: next_state = 3'b011;
        3'b011: begin
            done = 1'b1;
            out_bytes = {byte1, byte2, byte3};
            next_state = 3'b000;
        end
        default: next_state = 3'b000;
    endcase

    valid_byte1 = (state == 3'b001);
    valid_byte2 = (state == 3'b010);
    valid_byte3 = (state == 3'b011);
end

endmodule
