

module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

reg [4:0] state, next_state;
parameter WALK_LEFT = 5'b00001,
          WALK_RIGHT = 5'b00010,
          FALLING = 5'b00100,
          DIGGING = 5'b01000,
          SPLATTERED = 5'b10000;

reg [4:0] fall_counter;

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= WALK_LEFT;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        WALK_LEFT: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_right || dig)
                next_state = WALK_RIGHT;
            else
                next_state = WALK_LEFT;
        end
        
        WALK_RIGHT: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_left)
                next_state = WALK_LEFT;
            else
                next_state = WALK_RIGHT;
        end

        FALLING: begin
            if (fall_counter > 20 && ground) 
                next_state = SPLATTERED;
            else if (ground)
                next_state = state; // Continue in the same direction as before falling
            else
                next_state = FALLING;
        end
        
        DIGGING: begin
            if (!ground)
                next_state = FALLING;
            else if (bump_left || bump_right)
                next_state = state; // Continue digging, ignore bumps
            else
                next_state = state; // Continue digging until ground is 0
        end

        SPLATTERED: begin
            next_state = SPLATTERED;
        end
        
        default: 
            next_state = WALK_LEFT;
    endcase
end

always @(posedge clk or posedge areset) begin
    if (areset)
        fall_counter <= 0;
    else if (state == FALLING && !ground)
        fall_counter <= fall_counter + 1;
    else if (ground || state != FALLING)
        fall_counter <= 0;
end

assign walk_left = (state == WALK_LEFT);
assign walk_right = (state == WALK_RIGHT);
assign aaah = (state == FALLING) | (state == DIGGING && !ground);
assign digging = (state == DIGGING);

endmodule
