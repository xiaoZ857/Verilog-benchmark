
module TopModule (
  input a,
  input b,
  input cin,
  output cout,
  output sum
);


// VERILOG-EVAL: endmodule not found
