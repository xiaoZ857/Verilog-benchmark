
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  output walk_left,
  output walk_right,
  output aaah
);
always @(posedge clk or posedge areset) begin
    if (areset) begin
        walk_left <= 1'b1;
        walk_right <= 1'b0;
        aaah <= 1'b0;
    end else begin
        if (ground) begin
            aaah <= 1'b0;
            if (walk_left) begin
                if (bump_left) begin
                    walk_left <= 1'b0;
                    walk_right <= 1'b1;
                end else begin
                    walk_left <= 1'b1;
                    walk_right <= 1'b0;
                end
            end else if (walk_right) begin
                if (bump_right) begin
                    walk_left <= 1'b1;
                    walk_right <= 1'b0;
                end else begin
                    walk_left <= 1'b0;
                    walk_right <= 1'b1;
                end
            end
        end else begin
            aaah <= 1'b1;
        end
    end
end
endmodule
