
// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.
// The 7458 is a chip with four AND gates and two OR gates. Create a module
// in Verilog with the same functionality as the 7458 chip. It has 10 inputs
// and 2 outputs. You may choose to use an `assign` statement to drive each
// of the output wires, or you may choose to declare (four) wires for use as
// intermediate signals, where each internal wire is driven by the output of
// one of the AND gates.

module TopModule (
  input p1a,
  input p1b,
  input p1c,
  input p1d,
  input p1e,
  input p1f,
  output p1y,
  input p2a,
  input p2b,
  input p2c,
  input p2d,
  output p2y
);

// Implement p1y as the OR of two 3-input AND gates
assign p1y = (p1a & p1b & p1c) | (p1d & p1e & p1f);

// Implement p2y as the OR of two 2-input AND gates
assign p2y = (p2a & p2b) | (p2c & p2d);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
