
module TopModule (
  input c,
  input d,
  output [3:0] mux_in
);


// VERILOG-EVAL: endmodule not found
