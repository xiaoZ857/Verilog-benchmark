

module TopModule (
  output out
);

output out = 0;
endmodule
