
// TopModule.v
// -------------
// A module with no inputs and a single output that is permanently driven low.
// No clock or other logic is required.

`timescale 1ns / 1ps   // (optional – useful for simulation)

module TopModule (
    output out          // single output port
);

// Continuous assignment – drives the output low at all times
assign out = 1'b0;

endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
