
module TopModule (
  input c,
  input d,
  output [3:0] mux_in
);

// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.
// For the following Karnaugh map, give the circuit implementation using one
// 4-to-1 multiplexer and as many 2-to-1 multiplexers as required, but using
// as few as possible. You are not allowed to use any other logic gate and
// you must use _a_ and _b_ as the multiplexer selector inputs, as shown on
// the 4-to-1 multiplexer below.
//
//       ab
//   cd  00  01  11  10
//   00 | 0 | 0 | 0 | 1 |
//   01 | 1 | 0 | 0 | 0 |
//   11 | 1 | 0 | 1 | 1 |
//   10 | 1 | 0 | 0 | 1 |
//
// Consider a block diagram with inputs 'c' and 'd' going into a module
// called "top_module". This "top_module" has four outputs, mux_in[3:0],
// that connect to a four input mux. The mux takes as input {a,b} and ab =
// 00 is connected to mux_in[0], ab=01 is connected to mux_in[1], and so in.
// You are implementing in Verilog just the portion labelled "top_module",
// such that the entire circuit (including the 4-to-1 mux) implements the
// K

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
