
module TopModule (
  input [99:0] a,
  input [99:0] b,
  input sel,
  output [99:0] out
);
Here's the implementation of a 2:

// VERILOG-EVAL: endmodule not found
