
module TopModule (
  input clk,
  input d,
  output reg q
);
// Use two flip-flops: one triggered on positive edge, one on negative edge.
// Then combine their outputs with a multiplexer that toggles on the clock.
reg q_pos, q_neg;

always @(posedge clk) begin
    q_pos <= d;
end

always @(negedge clk) begin
    q_neg <= d;
end

always @(*) begin
    if (clk) begin
        q = q_pos;
    end else begin
        q = q_neg;
    end
end

endmodule
