

module TopModule (
  input clk,
  input reset,
  input [31:0] in,
  output reg [31:0] out
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        out <= 32'b0;
    end else begin
        for (int i = 0; i < 32; i++) begin
            if (in[i] == 1'b0 && out[i] == 1'b1) begin
                out[i] <= 1'b1;
            end else if (reset) begin
                out[i] <= 1'b0;
            end
        end
    end
end

always @(negedge clk or posedge reset) begin
    if (reset) begin
        // No action needed on negative edge for this logic
    end else begin
        for (int i = 0; i < 32; i++) begin
            if (in[i] == 1'b1 && out[i] == 1'b1) begin
                out[i] <= 1'b0;
            end
        end
    end
end

endmodule
