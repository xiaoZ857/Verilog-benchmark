

module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        q <= 32'h1;
    end else begin
        q[31:1] <= q[30:0];
        q[0] <= q[31] ^ q[21] ^ q[1] ^ q[0];
    end
end

endmodule
