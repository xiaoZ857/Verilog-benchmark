

module TopModule (
  input clock,
  input a,
  output reg p,
  output reg q
);

always @(posedge clock) begin
  if (a == 0) begin
    if (clock == 0) begin
      p <= 0;
      q <= 0;
    end else begin
      if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (clock == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <= 0;
        q <= 0;
      end else if (a == 0) begin
        p <=

// VERILOG-EVAL: endmodule not found
