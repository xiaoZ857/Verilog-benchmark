
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
  // State encoding (using binary encoding for clarity)
  parameter A = 3'b000,
            B = 3'b001,
            C = 3'b010,
            D = 3'b011,
            E = 3'b100,
            F = 3'b101;

  reg [2:0] current_state, next_state;

  // State register
  always @(posedge clk or posedge reset) begin
    if (reset)
      current_state <= A;
    else
      current_state <= next_state;
  end

  // Next state logic
  always @(*) begin
    case (current_state)
      A: next_state = (w == 1'b0) ? B : A;
      B: next_state = (w == 1'b0) ? C : D;
      C: next_state = (w == 1'b0) ? E : D;
      D: next_state = (w == 1'b0) ? F : A;
      E: next_state = (w == 1'b0) ? E : D;
      F: next_state = (w == 1'b0) ? C : D;
      default: next_state = A;
    endcase
  end

  // Output logic (Moore: output depends only on current_state)
  assign z = (current_state == E || current_state == F);

endmodule
