
module TopModule (
    input [5:0] y,
    input w,
    output Y1,
    output Y3
);

// State machine logic
assign Y1 = (y[4] == 0) && (y[5] == 0) ? w : (y[4] == 0) && (y[5] == 1) ? w : (y[2] == 0) && (y[3] == 0) ? w : (y[2] == 0) && (y[3] == 1) ? w : (y[1] == 0) && (y[3] == 0) ? w : (y[1] == 0) && (y[3] == 1) ? w : (y[4] == 1) && (y[5] == 0) ? w : (y[4] == 1) && (y[5] == 1) ? w;

assign Y3 = (y[4] == 0) && (y[5] == 0) ? w : (y[2] == 0) && (y[3] == 0) ? w : (y[1] == 0) && (y[3] == 0) ? w : (y[4] == 1) && (y[5] == 0) ? w : (y[2] == 1) && (y[3] == 0) ? w : (y[1] == 1) && (y[3] == 0) ? w : (y[4] == 1) && (y[5] == 1) ? w;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
