
module TopModule (
  input wire clk,
  input wire reset,
  input wire data,
  output wire [3:0] count,
  output reg counting,
  output reg done,
  input wire ack
);
always @(posedge clk) begin
    if (reset) begin
        counting <= 0;
        delay <= 4'b0;
        done <= 0;
        state = START;
    end

    case (state)
        START: begin
            if (data == 4'b1101) begin
                count <= data; // Store the start sequence pattern in count
                state = DELAY_SETUP;
            end
        end
        DELAY_SETUP: begin
            if (count[3] == 1 && count[2] == 1 && count[0] == 1) begin
                delay = count[1:0]; // Store the number of clock cycles to wait in delay
                state = COUNTING;
                counting <= 1;
            end
        end
        COUNTING: begin
            if (counting && rem_time > 0) begin
                rem_time--;
                if (rem_time == delay) begin
                    count <= delay; // Output the current remaining time
                end
                else begin
                    count <= rem_time + delay - 1; // Output the remaining time until timeout
                end
            end
            else if (counting && rem_time == 0) begin
                done <= 1; // Notify the user that the timer has timed out
                state = WAITING_ACK;
            end
        end
        WAITING_ACK: begin
            if (ack) begin
                count <= 4'bx; // Don't care value for count when waiting for ack
                state = START;
            end
        end
    endcase
end

// timescale directive outside the module definition
#timescale 1ns / 1ps
// default_nettype directives outside the module definitions
default_nettype register

// VERILOG-EVAL: endmodule not found
