

module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);



// VERILOG-EVAL: endmodule not found
