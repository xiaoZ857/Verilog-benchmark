

module TopModule (
  input clk,
  input reset,
  output shift_ena
);

  reg [1:0] state;
  reg shift_ena_reg;

  always @(posedge clk) begin
    if (reset) begin
      state <= 0;
      shift_ena_reg <= 1;
    end else begin
      case (state)
        0: begin
          shift_ena_reg <= 1;
          state <= 1;
        end
        1: begin
          shift_ena_reg <= 1;
          state <= 2;
        end
        2: begin
          shift_ena_reg <= 1;
          state <= 3;
        end
        3: begin
          shift_ena_reg <= 1;
          state <= 0;
        end
        default: begin
          state <= 0;
          shift_ena_reg <= 0;
        end
      endcase
    end
  end

  assign shift_ena = shift_ena_reg;
endmodule
