
module TopModule (
  output one
);
  
  // Assign the output to logic high (1)
  assign one = 1;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
