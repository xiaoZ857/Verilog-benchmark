
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);
always @(posedge clk) begin
    if (reset) begin
        done <= 1'b0;
        out_bytes <= 24'b0;
    end else begin
        done <= 1'b0;
        if (in[3]) begin
            out_bytes[23:16] <= in;
        end else if (out_bytes[23:16] != 8'b0) begin
            out_bytes[15:8] <= in;
        end else if (out_bytes[15:8] != 8'b0) begin
            out_bytes[7:0] <= in;
            done <= 1'b1;
        end
    end
end
endmodule
