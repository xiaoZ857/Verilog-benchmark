

module TopModule (
  input a,
  input b,
  output out
);

assign out = a nor b;
endmodule
