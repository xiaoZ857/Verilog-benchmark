
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);

reg current_state;

// State register with async reset and next state logic
always @(posed

// VERILOG-EVAL: endmodule not found
