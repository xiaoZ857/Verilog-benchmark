
module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);

always @(posedge clk) begin
  if (reset) begin
    q <= 4'd1;  // Reset to 1
  end else if (q == 4'd10) begin
    q <= 4'd1;  // After 10, go back to 1
  end else begin
    q <= q + 1;  // Increment counter
  end
end
endmodule
