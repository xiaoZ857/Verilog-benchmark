
time  a  b  c  d  q
0ns   0  0  0  0  1
5ns   0  0  0  0  1
10ns  0  0  0  0  1
15ns  0  0  0  0  1
20ns  0  0  0  1  0
25ns  0  0  1  0  0
30ns  0  0  1  1  1
35ns  0  1  0  0  0
40ns  0  1  0  1  1
45ns  0  1  1  0  1
50ns  0  1  1  1  0
55ns  1  0  0  0  0
60ns  1  0  0  1  1
65ns  1  0  1  0  1
70ns  1  0  1  1  0
75ns  1  1  0  0  1
80ns  1  1  0  1  0
85ns  1  1  1  0  0
90ns  1  1  1  1  1

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
