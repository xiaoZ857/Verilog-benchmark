
module TopModule (
  input clk,
  input resetn,
  input in,
  output out
);
  reg dff1, dff2, dff3, dff4;
  
  always @(posedge clk) begin
    if (!resetn) begin
      dff1 <= 1'b0;
      dff2 <= 1'b0;
      dff3 <= 1'b0;
      dff4 <= 1'b0;
    end else begin
      dff1 <= in;
      dff2 <= dff1;
      dff3 <= dff2;
      dff4 <= dff3;
    end
  end
  
  assign out = dff4;
endmodule

// VERILOG-EVAL: errant inclusion of module definition
