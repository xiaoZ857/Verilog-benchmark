
// This timescale directive should be placed at the top of the file, not inside a module
`timescale 1ns / 1ps

module TopModule (
  input in1,
  input in2,
  input in3,
  output logic out
);

  // XNOR and XOR implementation
  wire xnor_out;
  
  // XNOR gate: (in1 == in2) is equivalent to !XOR
  assign xnor_out = (in1 == in2);
  
  // XOR gate with second input in3
  assign out = xnor_out ^ in3;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
