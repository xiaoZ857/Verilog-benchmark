
module TopModule (
  input [4:1] x,
  output logic f
);
assign f = (~x[3] & x[4] & x[2] & x[1]) |  // x[3]x[4]=01, x[1]x[2]=11
           (x[3] & ~x[4] & ~x[2]) |        // x[3]x[4]=10, x[1]x[2]=00,01 (both 1)
           (x[3] & ~x[4] & x[1]) |         // x[3]x[4]=10, x[1]x[2]=01,11
           (x[3] & x[4] & ~x[1]) |         // x[3]x[4]=11, x[1]x[2]=00,10
           (x[3] & x[4] & ~x[2]);          // x[3]x[4]=11, x[1]x[2]=00,01
