
module TopModule (
  input [5:0] y,
  input w,
  output Y1,
  output Y3
);
  // Y1 is the input to the flip-flop for state y[1] (B)
  // From the state diagram:
  //  - If in state A (000001), on input 0, stay in A.  Y1 = 0
  //  - If in state A (000001), on input 1, go to B.  Y1 = 1
  //  - If in state B (000010), on input 0, go to D.  Y1 = 0
  //  - If in state B (000010), on input 1, go to C.  Y1 = 1
  always_comb begin
    if (y == 6'b000001) begin // State A
      Y1 = w;
    end else if (y == 6'b000010) begin // State B
      Y1 = w;
    end else begin
      Y1 = 1'b0; // Default: stay in current state (not strictly needed)
    end
  end

  // Y3 is the input to the flip-flop for state y[3] (D)
  // From the state diagram:
  //  - If in state A (000001), on input 0, stay in A.  Y3 = 0
  //  - If in state A (000001), on input 1, go to B.  Y3 = 0
  //  - If in state B (000010), on input 0, go to D.  Y3 = 0
  //  - If in state B (000010), on input 1, go to C.  Y3 = 0
  //  - If in state C (000100), on input 0, go to D.  Y3 = 0
  //  - If in state C (000100), on input 1, go to E.  Y3 = 1
  //  - If in state D (001000), on input 0, go to A.  Y3 = 0
  //  - If in state D (001000), on input 1, go to F.  Y3 = 1
  //  - If in state E (010000), on input 0, go to D.  Y3 = 0
  //  - If in state E (010000), on input 1, go to E.  Y3 = 1
  //  - If in state F (100000), on input 0, go to D.  Y3 = 0
  //  - If in state F (100000), on input 1, go to C.  Y3 = 1
  always_comb begin
    if (y == 6'b000001) begin // State A
      Y3 = 1'b0;
    end else if (y == 6'b000010) begin // State B
      Y3 = 1'b0;
    end else if (y == 6'b000100) begin // State C
      Y3 = w;
    end else if (y == 6'b001000) begin // State D
      Y3 = w;
    end else if (y == 6'b010000) begin // State E
      Y3 = w;
    end else if (y == 6'b100000) begin // State F
      Y3 = w;
    end else begin
      Y3 = 1'b0; // Default: stay in current state (not strictly needed)
    end
  end

endmodule
