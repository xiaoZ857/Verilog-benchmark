

module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);

module FSMDatapath (
  input clk,
  input [7:0] in,
  input reset,
  output reg [23:0] out_bytes,
  output reg done
);

reg [2:0] state; // State machine registers
always @(posedge clk) begin
  if (reset) begin
    state <= 4'b0001; // Reset to initial state
  end else begin
    case (state)
      4'b0001: begin // Idle state
        if (in[3] == 1) state <= 4'b0010; // Transition to message receiving state when in[3]=1
      end
      4'b0010: begin // Message receiving state
        out_bytes <= in; // Store the received byte in out_bytes
        if (out_bytes == 24'h0000_0000_0000_0009) state <= 4'b0100; // Transition to done state when message is complete
        else state <= 4'b0010; // Stay in message receiving state if message is not complete
      end
      4'b0100: begin // Done state
        out_bytes <= {out_bytes[23:16], out_bytes[15:8], out_bytes[7:0]}; // Reorder the bytes in out_bytes
        done <= 1'b1; // Signal that a message has been received
        state <= 4'b1000; // Transition to idle state after signaling done
      end
      4'b1000: begin // Idle state
        done <= 1'b0; // Reset done signal
      end
    endcase
  end
end

// Add any necessary initializations and testbench code here

endmodule
