
module TopModule (
  input [4:0] a,
  input [4:0] b,
  input [4:0] c,
  input [4:0] d,
  input [4:0] e,
  input [4:0] f,
  output [7:0] w,
  output [7:0] x,
  output [7:0] y,
  output [7:0] z
);
assign w = {a, b, c, d, e, f, 1'b0, 1'b0};
assign x = {f, e, d, c, b, a, 1'b0, 1'b0};
assign y = {c, b, a, f, e, d, 1'b0, 1'b0};
assign z = {d, e, f, g, h, i, j, k};

// VERILOG-EVAL: endmodule not found
