
module TopModule (
  output out
);

  // Assign logic low (0) to the output
  assign out = 1'b0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
