
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);
WALK_L, WALK_R, FALL_L, FALL_R, DIG_L, DIG_R, SPLATTER

// VERILOG-EVAL: abnormal backticks count
