
// ------------------------------------------------------------
//  2‑to‑1 Multiplexer (100‑bit wide)
//  When sel = 0 → out = a
//  When sel = 1 → out = b
// ------------------------------------------------------------
`timescale 1ns / 1ps

module TopModule (
    input  wire [99:0] a,   // First 100‑bit input
    input  wire [99:0] b,   // Second 100‑bit input
    input  wire        sel, // Select signal
    output wire [99:0] out  // 100‑bit output
);

    // Combinational assignment – synthesizable
    assign out = sel ? b : a;

    // Alternative (always @* block) – equivalent
    // always @* begin
    //     if (sel)
    //         out = b;
    //     else
    //         out = a;
    // end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
