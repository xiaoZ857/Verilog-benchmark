
module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);
always @(posedge clk or posedge reset) begin
    if (reset) begin
        q <= 4'b0000; // Synchronous active-high reset
    end else begin
        if (q == 4'b1111) begin
            q <= 4'b0000; // Wrap around to 0 when it reaches 15
        end else begin
            q <= q + 1;   // Regular increment otherwise
        end
    end
end

endmodule
