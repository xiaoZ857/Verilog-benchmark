
module TopModule (
  input [1023:0] in,
  input [7:0] sel,
  output [3:0] out
);
  // Calculate the starting index of the selected input based on the selector.
  wire [9:0] index;
  assign index = sel * 4;

  // Select the 4-bit input based on the calculated index.
  assign out = in[index + 3 : index];

endmodule
