
assign f = x[1]'x[2] & x[3]' | x[1]'x[4];

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
