
module TopModule (
    input clk,
    input load,
    input ena,
    input [1:0] amount,
    input [63:0] data,
    output reg [63:0] q
);

    always @(posedge clk) begin
        if (load) begin
            // Load the data into the register when load is active high
            q <= data;
        end else if (ena) begin
            case (amount)
                2'b00: begin
                    // Shift left by 1 bit
                    q <= {q[62:0], 1'b0};
                end
                2'b01: begin
                    // Shift left by 8 bits
                    q <= {q[55:0], 8'b00000000};
                end
                2'b10: begin
                    // Arithmetic right shift by 1 bit (sign extension)
                    q <= {q[63], q[62:0]};
                end
                2'b11: begin
                    // Arithmetic right shift by 8 bits (sign extension)
                    q <= {q[63:56], q[55:0]};
                end
            endcase
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
