
module TopModule (
  input in,
  output out
);
 ```verilog
assign out = in;
endmodule

// VERILOG-EVAL: abnormal backticks count
