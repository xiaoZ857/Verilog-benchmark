
module TopModule (
    input  wire clk,    // clock
    input  wire j,      // input that drives OFF →

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
