
module TopModule (
  input clk,
  input reset,
  input ena,
  output reg pm,
  output reg [7:0] hh,
  output reg [7:0] mm,
  output reg [7:0] ss
);
assign pm = (reset || ena) ? 1'b0 : (clk == 1'b1);
always @(posedge clk) begin
    if (ena)
        hh <= {hh[1], hh[0] + 1};
    else if (reset)
        hh <= 7'b00000;
end

assign mm = (hh[1] == 1'b1) ? 7'b59 : hh[1:2];
assign ss = (mm[1] == 1'b1) ? 7'b59 : mm[1:2];

always @(posedge clk) begin
    if (ena)
        mm <= {mm[1], mm[0] + 1};
    else if (reset)
        mm <= 7'b00000;
end

assign ss = (mm[1] == 1'b1) ? 7'b59 : mm[1:2];

always @(posedge clk) begin
    if (ena)
        ss <= {ss[1], ss[0] + 1};
    else if (reset)
        ss <= 7'b00000;
end

assign hh = ((mm[1] == 1'b1) ? mm : mm[1:2]) * 10 + hh[1];

endmodule
