
// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.

// Moore state machine with two states, two inputs, and one output.
// Reset is an active-high asynchronous reset to state OFF.

module TopModule (
  input clk,
  input j,
  input k,
  input areset,
  output out
);

  reg [1:0] state;
  
  always @(posedge clk or posedge areset) begin
    if (areset) begin
      state <= 2'b00; // OFF state
    end else case (state)
      2'b00: begin // OFF state
        if (j == 1) state <= 2'b01; // ON state
        else state <= 2'b00;
      end
      2'b01: begin // ON state
        if (k == 1) state <= 2'b00; // OFF state
        else state <= 2'b01;
      end
    endcase
  end

  assign out = (state == 2'b01) ? 1 : 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
