
module TopModule (
  input clk,
  input reset,
  input x,
  output reg z
);
always @(posedge clk) begin
    if (reset)
        {q2, q1, q0} <= 3'b000;
    else begin
        case ({q2, q1, q0})
            3'b000: 
                if (x == 0) {q2, q1, q0} <= 3'b000; else {q2, q1, q0} <= 3'b001;
                z = 0;
            3'b001: 
                if (x == 0) {q2, q1, q0} <= 3'b001; else {q2, q1, q0} <= 3'b100;
                z = 0;
            3'b010: 
                if (x == 0) {q2, q1, q0} <= 3'b010; else {q2, q1, q0} <= 3'b001;
                z = 0;
            3'b011: 
                if (x == 0) {q2, q1, q0} <= 3'b010; else {q2, q1, q0} <= 3'b011;
                z = 1;
            3'b100: 
                if (x == 0) {q2, q1, q0} <= 3'b011; else {q2, q1, q0} <= 3'b100;
                z = 1;
            default: 
                {q2, q1, q0} <= {q2, q1, q0};
        endcase
    end
end

endmodule
