
`timescale 1ns / 1ps

module TopModule (
    input  wire        clk,   // clock input
    input  wire        reset, // active‑high synchronous reset
    output reg  [3:0]  q     // 4‑bit counter output
);

    // Synchronous logic: triggered on the rising edge of clk
    always @(posedge clk) begin
        if (reset) begin
            // Reset is synchronous – performed on the clock edge
            q <= 4'd0;
        end
        else begin
            // Count from 0 to 9, then wrap to 0
            if (q == 4'd9) begin
                q <= 4'd0;
            end
            else begin
                q <= q + 1'b1;
            end
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
