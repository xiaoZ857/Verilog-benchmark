
module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);
reg state;
reg next_state;

always @(*) begin
    case (state)
        1'b0: next_state = j ? 1'b1 : 1'b0;
        1'b1: next_state = k ? 1'b0 : 1'b1;
        default: next_state = 1'b0;
    endcase
end

always @(posedge clk) begin
    if (reset)
        state <= 1'b0;
    else
        state <= next_state;
end

assign out = state;
endmodule
