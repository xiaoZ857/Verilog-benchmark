
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output reg walk_left = 1'b0,
  output reg walk_right = 1'b0,
  output reg aaah = 1'b0,
  output reg digging = 1'b0
);

    // Define states
    typedef enum logic [2:0] {
        WALK_LEFT,       // Lemming walks left
        WALK_RIGHT,      // Lemming walks right
        FALLING,         // Lemming is falling and saying "aaah!"
        DIGGING          // Lemming is digging
    } state_t;

    state_t current_state, next_state;

    always_ff @(posedge clk or posedge areset) begin
        if (areset)
            current_state <= WALK_LEFT; // Asynchronous reset to walk left
        else
            current_state <= next_state;
    end

    always_comb begin
        // Default outputs for each state transition
        walk_left = 1'b0;
        walk_right = 1'b0;
        aaah = 1'b0;
        digging = 1'b0;

        case (current_state)
            WALK_LEFT: begin
                if (!ground) begin
                    next_state = FALLING; // Fall when ground disappears
                    aaah = 1'b1;
                end else if (bump_right || dig) begin
                    next_state = (dig) ? DIGGING : WALK_RIGHT; // Dig or switch to walking right
                    digging = (dig) ? 1'b1 : 1'b0;
                end else if (bump_left) begin
                    next_state = WALK_LEFT; // Remain walking left when bumped on the left only
                end else begin
                    next_state = WALK_LEFT; // Continue walking left
                    walk_left = 1'b1;
                end
            end

            WALK_RIGHT: begin
                if (!ground) begin
                    next_state = FALLING;
                    aaah = 1'b1;
                end else if (bump_left || dig) begin
                    next_state = (dig) ? DIGGING : WALK_LEFT; // Dig or switch to walking left
                    digging = (dig) ? 1'b1 : 1'b0;
                end else if (bump_right) begin
                    next_state = WALK_RIGHT; // Remain walking right when bumped on the right only
                end else begin
                    next_state = WALK_RIGHT; // Continue walking right
                    walk_right = 1'b1;
                end
            end

            FALLING: begin
                if (ground) begin
                    next_state = current_state == WALK_LEFT ? WALK_LEFT : WALK_RIGHT; // Resume previous direction
                end else begin
                    next_state = FALLING; // Continue falling
                    aaah = 1'b1;
                end
            end

            DIGGING: begin
                if (!ground) begin
                    next_state = FALLING;
                    aaah = 1'b1;
                end else begin
                    next_state = current_state == WALK_LEFT ? WALK_LEFT : WALK_RIGHT; // Resume previous direction when ground appears
                    digging = 1'b1;
                end
            end

        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
