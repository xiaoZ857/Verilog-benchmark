

module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] pedge
);



// VERILOG-EVAL: endmodule not found
