

module TopModule (
  input in,
  input [3:0] state,
  output reg [3:0] next_state,
  output out
);

  always @(in, state) begin
    case (state)
      4'b0001: begin // State A
        if (in == 0)
          next_state = 4'b0001;
        else
          next_state = 4'b0010;
        out = 0;
      end
      4'b0010: begin // State B
        if (in == 0)
          next_state = 4'b0100;
        else
          next_state = 4'b0010;
        out = 0;
      end
      4'b0100: begin // State C
        if (in == 0)
          next_state = 4'b0001;
        else
          next_state = 4'b1000;
        out = 0;
      end
      4'b1000: begin // State D
        if (in == 0)
          next_state = 4'b0100;
        else
          next_state = 4'b0010;
        out = 1;
      end
    endcase
  end

endmodule
