
module TopModule (
  input clk,
  input d,
  input ar,
  output logic q
);


// VERILOG-EVAL: endmodule not found
