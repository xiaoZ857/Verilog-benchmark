

module TopModule (
  input clk,
  input areset,
  input train_valid,
  input train_taken,
  output logic [1:0] state
);



// VERILOG-EVAL: endmodule not found
