
// Define the module TopModule that implements the Game of Life
module TopModule (
  // Clock and load signals
  input clk,
  input load,
  
  // Data for loading initial state
  input [255:0] data,
  
  // Output vector representing the current game state
  output reg [255:0] q
);

// Initialize signal to store the previous game state (for calculating neighbors)
reg [255:0] prev_q;

// Calculate the number of neighbors for each cell in the grid
always_ff @(posedge clk) begin
  // Store the current state in prev_q before changing it
  prev_q <= q;
  
  // Iterate over each cell in the grid (16x16)
  for (int i = 0; i < 256; i++) begin
    int j = (i % 16); // Calculate row and column indices
    
    // Initialize variables to store the number of live neighbors
    int live_neighbors = 0;
    
    // Iterate over each neighbor in a toroid boundary around cell (i, j)
    for (int x = -1; x <= 1; x++) begin
      for (int y = -1; y <= 1; y++) begin
        if ((x == 0) && (y == 0)) continue;
        
        int neighbor_i = i + x * 16;
        int neighbor_j = j + y;
        
        // Calculate the toroid boundary condition to wrap around
        neighbor_i %= 256;
        neighbor_j %= 16;
        
        if (prev_q[neighbor_i + neighbor_j * 16] == 1) begin
          live_neighbors++;
        end
      end
    end
    
    // Apply the Game of Life rules based on the number of neighbors
    q[i] = (live_neighbors == 0) ? 0 : ((live_neighbors == 2) || (live_neighbors == 3)) ? q[i] : 1;
  end
end

// Load initial state from data on rising edge of load signal
always_ff @(posedge load) begin
  q <= data;
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
