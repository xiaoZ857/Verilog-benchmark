
`timescale 1ns / 1ps

module TopModule (
    input  [99:0] in,
    output reg [99:0] out
);

    /*------------------------------------------------------------
     *  Reverse the bit order of the 100‑bit input vector.
     *  out[0]  = in[99]
     *  out[1]  = in[98]
     *  ...
     *  out[99] = in[0]
     *------------------------------------------------------------*/
    always @(*) begin
        integer i;
        for (i = 0; i < 100; i = i + 1) begin
            out[i] = in[99 - i];
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
