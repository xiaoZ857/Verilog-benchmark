
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
  // State encoding: A=00, B=01, C=10, D=11
  reg [1:0] state, next_state;
  
  // State register with synchronous reset
  always @(posedge clk) begin
    if (reset)
      state <= 2'b00; // Reset to state A
    else
      state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      2'b00: // State A
        next_state = in ? 2'b01 : 2'b00; // A->B if in=1, else stay A
      2'b01: // State B
        next_state = in ? 2'b01 : 2'b10; // B->C if in=0, else stay B
      2'b10: // State C
        next_state = in ? 2'b11 : 2'b00; // C->D if in=1, else go to A
      2'b11: // State D
        next_state = in ? 2'b01 : 2'b10; // D->B if in=1, else go to C
      default:
        next_state = 2'b00; // Default to state A
    endcase
  end
  
  // Output logic (Moore: output depends only on state)
  assign out = (state == 2'b11); // Output 1 only in state D

endmodule
