
module TopModule (
  input d,
  input done_counting,
  input ack,
  input [9:0] state, // 10-bit one-hot current state
  output B3_next,
  output S_next,
  output S1_next,
  output Count_next,
  output Wait_next,
  output done,
  output counting,
  output shift_ena
);

  // Next state logic
  assign B3_next = state[6]; // From B2 state
  assign S_next = (state[0] & ~d) | (state[1] & ~d) | (state[3] & ~d) | (state[9] & ack); // From S(d=0), S1(d=0), S110(d=0), Wait(ack=1)
  assign S1_next = state[0] & d; // From S state with d=1
  assign Count_next = state[7] | (state[8] & ~done_counting); // From B3 state or Count state with done_counting=0
  assign Wait_next = (state[8] & done_counting) | (state[9] & ~ack); // From Count state with done_counting=1 or Wait state with ack=0
  
  // Output logic
  assign shift_ena = state[4] | state[5] | state[6] | state[7]; // Active in B0, B1, B2, B3 states
  assign counting = state[8]; // Active in Count state
  assign done = state[9]; // Active in Wait state
endmodule
