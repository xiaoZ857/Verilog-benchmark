

module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);



// VERILOG-EVAL: endmodule not found
