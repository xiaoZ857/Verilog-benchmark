
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);

reg [2:0] current_state, next_state;

// State encoding
parameter A = 3'b000;
parameter B = 3'b001;
parameter C = 3'b010;
parameter D = 3'b011;
parameter E = 3'b100;
parameter F = 3'b101;

// State transition logic
always @(posedge clk) begin
  if (reset) begin
    current_state <= A;
  end else begin
    current_state <= next_state;
  end
end

// Next state logic
always @(*) begin
  case (current_state)
    A: begin
      if (w) next_state = A;
      else next_state = B;
    end
    B: begin
      if (w) next_state = D;
      else next_state = C;
    end
    C: begin
      if (w) next_state = D;
      else next_state = E;
    end
    D: begin
      if (w) next_state = A;
      else next_state = F;
    end
    E: begin
      if (w) next_state = D;
      else next_state = E;
    end
    F: begin
      if (w) next_state = D;
      else next_state = C;
    end
    default: next_state = A;
  endcase
end

// Output logic
always @(*) begin
  case (current_state)
    E: z = 1'b1;
    F: z = 1'b1;
    default: z = 1'b0;
  endcase
end

endmodule
