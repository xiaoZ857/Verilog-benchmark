
module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);
always @(posedge clk or negedge aresetn) begin
    if (!aresetn) begin
        z <= 0; // Reset output to logic-0 when asynchronous reset is asserted
    end else begin
        case (current_state)
            IDLE:
                if (x == 1'b1) begin
                    current_state = WAIT_FOR_ONE;
                end
                break;
            WAIT_FOR_ONE:
                if (x == 1'b0) begin
                    current_state = WAIT_FOR_TWO;
                end else begin
                    z <= 0; // Reset output to logic-0 when first '1' is followed by '0'
                    current_state = IDLE;
                end
                break;
            WAIT_FOR_TWO:
                if (x == 1'b1) begin
                    z <= 1; // Assert output to logic-1 when second '0' is followed by '1'
                    current_state = IDLE;
                end else begin
                    z <= 0; // Reset output to logic-0 when second '0' is not followed by '1'
                    current_state = IDLE;
                end
        endcase
    end
end

endmodule
