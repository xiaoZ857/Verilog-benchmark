
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

reg [2:0] state, next_state;
reg [4:0] fall_counter;
reg walking_left; // Track current walking direction

parameter WALK_LEFT = 3'b000;
parameter WALK_RIGHT = 3'b001;
parameter FALLING = 3'b010;
parameter DIGGING = 3'b011;
parameter SPLATTERED = 3'b100;

always @(posedge clk or posedge areset) begin
  if (areset) begin
    state <= WALK_LEFT;
    fall_counter <= 5'b0;
    walking_left <= 1'b1; // Start walking left
  end else begin
    state <= next_state;
    if (state == FALLING) begin
      fall_counter <= fall_counter + 1;
    end else begin
      fall_counter <= 5'b0;
    end
    // Update walking direction when switching between WALK_LEFT and WALK_RIGHT
    if (next_state == WALK_LEFT) begin
      walking_left <= 1'b1;
    end else if (next_state == WALK_RIGHT) begin
      walking_left <= 1'b0;
    end
  end
end

always @(*) begin
  next_state = state;
  case (state)
    WALK_LEFT: begin
      // Priority: fall > dig > switch directions
      if (!ground) begin
        next_state = FALLING;
      end else if (dig) begin
        next_state = DIGGING;
      end else if (bump_left || bump_right) begin
        next_state = WALK_RIGHT;
      end
    end
    
    WALK_RIGHT: begin
      // Priority: fall > dig > switch directions
      if (!ground) begin
        next_state = FALLING;
      end else if (dig) begin
        next_state = DIGGING;
      end else if (bump_left || bump_right) begin
        next_state = WALK_LEFT;
      end
    end
    
    FALLING: begin
      if (

// VERILOG-EVAL: endmodule not found
