
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);

  always @(posedge clk) begin
    case (y[3:1])
      4'0000: Y2 <= 0; // A (0) --0--> B, A (0) --1--> A
      4'0001: Y2 <= 0; // B (0) --0--> C, B (0) --1--> D
      4'0010: Y2 <= 0; // C (0) --0--> E, C (0) --1--> D
      4'0011: Y2 <= 0; // D (0) --0--> F, D (0) --1--> A
      4'0100: Y2 <= 0; // E (1) --0--> E, E (1) --1--> D
      4'0101: Y2 <= 0; // F (1) --0--> C, F (1) --1--> D
      default: Y2 <= 0;
    endcase
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
