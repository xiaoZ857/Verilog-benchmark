
module TopModule (
  input [7:0] in,
  output [31:0] out
);
wire signed [7:0] sign_in; // Extract the sign bit from the input
assign sign_in = in[7];

// Create a 24-bit constant for replication
parameter sign_repl [23:0] = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                               1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                               1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};

// Replicate the sign bit and concatenate with the input
wire [31:0] temp_out;
for(int i = 0; i < 24; i++)
    temp_out[i + 8] = sign_repl[i];
temp_out[8:0] = in;

assign out = temp_out; // Assign the result to output

endmodule
