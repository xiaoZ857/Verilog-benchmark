
module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);

always @(posedge clk) begin
  if (load) begin
    q <= data;
  end else begin
    integer i, j, neighbor_count;
    reg [255:0] next_q;
    
    next_q = 256'b0;
    
    for (i = 0; i < 16; i = i + 1) begin
      for (j = 0; j < 16; j = j + 1) begin
        neighbor_count = 0;
        
        // Calculate neighbors with toroidal wrapping
        // Top row neighbors
        neighbor_count = neighbor_count + q[((i+15)%16)*16 + ((j+15)%16)];
        neighbor_count = neighbor_count + q[((i+15)%16)*16 + j];
        neighbor_count = neighbor_count + q[((i+15)%16)*16 + ((j+1)%16)];
        
        // Middle row neighbors
        neighbor_count = neighbor_count + q[i*16 + ((j+15)%16)];
        neighbor_count = neighbor_count + q[i*16 + ((j+1)%16)];
        
        // Bottom row neighbors
        neighbor_count = neighbor_count + q[((i+1)%16)*16 + ((j+15)%16)];
        neighbor_count = neighbor_count + q[((i+1)%16)*16 + j];
        neighbor_count = neighbor_count + q[((i+1)%16)*16 + ((j+1)%16)];
        
        // Apply Game of Life rules
        if (neighbor_count <= 1) begin
          next_q[i*16 + j] = 1'b0;
        end else if (neighbor_count == 2) begin
          next_q[i*16 + j] = q[i*16 + j];
        end else if (neighbor_count == 3) begin
          next_q[i*16 + j] = 1'b1;
        end else begin
          next_q[i*16 + j] = 1'b0;
        end
      end
    end
    
    q <= next_q;
  end
end
endmodule
