
module TopModule (
  input clk,
  input a,
  output reg q
);
always @(posedge clk) begin
    if (a == 1 && q == 0) begin
        q <= 1;
    end else if (a == 0 && q == 1) begin
        q <= 0;
    end else if (a == 1 && q == 1) begin
        q <= q; // Keep the current state
    end else if (a == 0 && q == 0) begin
        q <= 0;
    end
end

// VERILOG-EVAL: endmodule not found
