
// TopModule.v
// 10‑bit synchronous counter that counts from 0 to 999 inclusive.
// The counter wraps back to 0 after reaching 999 (period = 1000 cycles).
// `reset` is active‑high and synchronous.

`timescale 1ns / 1ps

module TopModule (
    input  wire        clk,   // Positive‑edge clock
    input  wire        reset, // Active‑high synchronous reset
    output reg  [9:0]  q      // 10‑bit counter output
);

    // --------------------------------------------------------------------
    // Parameters
    // --------------------------------------------------------------------
    localparam MAX_COUNT = 10'd999;   // Final count value (0‑999)

    // --------------------------------------------------------------------
    // Counter logic
    // --------------------------------------------------------------------
    always @(posedge clk) begin
        if (reset) begin
            q <= 10'd0;               // Reset to zero
        end
        else if (q == MAX_COUNT) begin
            q <= 10'd0;               // Wrap after reaching 999
        end
        else begin
            q <= q + 1'b1;            // Increment normally
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
