
module TopModule (
  input in,
  output out
);
  
  // Implement NOT gate using the NOT keyword
  assign out = !in;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
