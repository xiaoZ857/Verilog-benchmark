
module TopModule (
  input cpu_overheated,
  output reg shut_off_computer,
  input arrived,
  input gas_tank_empty,
  output reg keep_driving
);
module top_module (
    input      cpu_overheated,
    output reg shut_off_computer,
    input      arrived,
    input      gas_tank_empty,
    output reg keep_driving  
);

    always @(*) begin
        // Default assignments to prevent latches
        shut_off_computer = 0;
        
        if (cpu_overheated) begin
            shut_off_computer = 1;
        end
    end

    always @(*) begin
        // Default assignment to prevent latches
        keep_driving = 0;  // default value when arrived or gas_tank_empty
        
        if (~arrived && ~gas_tank_empty) begin
            keep_driving = 1;
        end
    end

endmodule
