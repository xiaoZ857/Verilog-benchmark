
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output q
);

assign q = (!a && !b && !c) || (!a && !b && d) || (!a && c && !d) || (!a && c && d) || (a && !b && !c) || (a && !b && d) || (a && c && !d) || (a && c && d) || (b && !c && !d) || (b && !c && d) || (b && c && !d) || (b && c && d) || (c && !d && !a) || (c && !d && a) || (c && d && !a) || (c && d && a);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
