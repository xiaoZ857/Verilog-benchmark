
module TopModule (
  input wire clk,
  input wire in,
  input wire reset,
  output reg out
);

  // State encoding
  typedef enum logic [1:0] {
    STATE_A = 2'b00,
    STATE_B = 2'b01,
    STATE_C = 2'b10,
    STATE_D = 2'b11
  } state_t;

  // Registers for current and next states
  state_t current_state, next_state;

  // Output logic based on the current state
  always @(*) begin
    case (current_state)
      STATE_A: out = 1'b0;
      STATE_B: out = 1'b0;
      STATE_C: out = 1'b0;
      STATE_D: out = 1'b1;
      default: out = 1'bx; // Undefined state
    endcase
  end

  // Next state logic
  always @(*) begin
    case (current_state)
      STATE_A: next_state = in ? STATE_B : STATE_A;
      STATE_B: next_state = in ? STATE_B : STATE_C;
      STATE_C: next_state = in ? STATE_D : STATE_A;
      STATE_D: next_state = in ? STATE_B : STATE_C;
      default: next_state = STATE_A; // Undefined state
    endcase
  end

  // State transition and reset logic
  always @(posedge clk or posedge reset) begin
    if (reset)
      current_state <= STATE_A;
    else
      current_state <= next_state;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
