
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);

// FSM for serial data reception with start/stop bits
reg [3:0] state, next_state;
reg [7:0] data_reg;
reg [2:0] bit_count;

// State definitions
localparam IDLE = 4'd0;
localparam START = 4'd1;
localparam DATA0 = 4'd2;
localparam DATA1 = 4'd3;
localparam DATA2 = 4'd4;
localparam DATA3 = 4'd5;
localparam DATA4 = 4'd6;
localparam DATA5 = 4'd7;
localparam DATA6 = 4'd8;
localparam DATA7 = 4'd9;
localparam STOP = 4'd10;
localparam WAIT_STOP = 4'd11;

// State register
always @(posedge clk) begin
    if (reset) begin
        state <= IDLE;
        data_reg <= 8'b0;
        bit_count <= 3'b0;
    end else begin
        state <= next_state;
        case (state)
            START: begin
                data_reg <= 8'b0;
                bit_count <= 3'b0;
            end
            DATA0, DATA1, DATA2, DATA3, DATA4, DATA5, DATA6: begin
                data_reg <= {in, data_reg[7:1]};
                bit_count <= bit_count + 1;
            end
            DATA7: begin
                data_reg <= {in, data_reg[7:1]};
            end
        endcase
    end
end

// Next state logic
always @(*) begin
    next_state = state;
    case (state)
        IDLE: begin
            if (in == 0) begin
                next_state = START;
            end
        end
        START: begin
            next_state = DATA0;
        end
        DATA0: next_state = DATA1;
        DATA1: next_state = DATA2;
        DATA2: next_state = DATA3;
        DATA3: next_state = DATA4;
        DATA4: next_state = DATA5;
        DATA5: next_state = DATA6;
        DATA6: next_state = DATA7;
        DATA7: next_state = STOP;
        STOP: begin
            if (in == 1) begin
                next_state = IDLE;
            end else begin
                next_state = WAIT_STOP;
            end
        end
        WAIT_STOP: begin
            if (in == 1) begin
                next_state = IDLE;
            end
        end
    endcase
end

// Output logic
assign out_byte = data_reg;
assign done = (state == STOP && in == 1);

endmodule
