
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

  reg [2:0] state, next_state;
  
  // State encoding
  localparam WALK_LEFT  = 3'b000;
  localparam WALK_RIGHT = 3'b001;
  localparam FALL_LEFT  = 3'b010;
  localparam FALL_RIGHT = 3'b011;
  localparam DIG_LEFT   = 3'b100;
  localparam DIG_RIGHT  = 3'b101;
  
  // State transition logic
  always @(*) begin
    case (state)
      WALK_LEFT: begin
        if (!ground) 
          next_state = FALL_LEFT;
        else if (dig) 
          next_state = DIG_LEFT;
        else if (bump_left || (bump_left && bump_right)) 
          next_state = WALK_RIGHT;
        else 
          next_state = WALK_LEFT;
      end
      
      WALK_RIGHT: begin
        if (!ground) 
          next_state = FALL_RIGHT;
        else if (dig) 
          next_state = DIG_RIGHT;
        else if (bump_right || (bump_left && bump_right)) 
          next_state = WALK_LEFT;
        else 
          next_state = WALK_RIGHT;
      end
      
      FALL_LEFT: begin
        if (ground) 
          next_state = WALK_LEFT;
        else 
          next_state = FALL_LEFT;
      end
      
      FALL_RIGHT: begin
        if (ground) 
          next_state = WALK_RIGHT;
        else 
          next_state = FALL_RIGHT;
      end
      
      DIG_LEFT: begin
        if (!ground) 
          next_state = FALL_LEFT;
        else 
          next_state = DIG_LEFT;
      end
      
      DIG_RIGHT: begin
        if (!ground) 
          next_state = FALL_RIGHT;
        else 
          next_state = DIG_RIGHT;
      end
      
      default: 
        next_state = WALK_LEFT;
    endcase
  end
  
  // State register
  always @(posedge clk or posedge areset) begin
    if (areset) 
      state <= WALK_LEFT;
    else 
      state <= next_state;
  end
  
  // Output logic (Moore machine)
  assign walk_left = (state == WALK_LEFT);
  assign walk_right = (state == WALK

// VERILOG-EVAL: endmodule not found
