
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
reg state;
reg next_state;

always @(posedge clk) begin
    if (reset)
        state <= 1'b0;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        1'b0: next_state = in ? 1'b0 : 1'b1;
        1'b1: next_state = in ? 1'b1 : 1'b0;
        default: next_state = 1'b0;
    endcase
end

assign out = (state == 1'b0) ? 1'b1 : 1'b0;

endmodule
