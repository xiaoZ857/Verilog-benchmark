
module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] pedge
);
assign pedge[0] = (in[0] == 0) && (in[0] != 0);
assign pedge[1] = (in[1] == 0) && (in[1] != 0);
assign pedge[2] = (in[2] == 0) && (in[2] != 0);
assign pedge[3] = (in[3] == 0) && (in[3] != 0);
assign pedge[4] = (in[4] == 0) && (in[4] != 0);
assign pedge[5] = (in[5] == 0) && (in[5] != 0);
assign pedge[6] = (in[6] == 0) && (in[6] != 0);
assign pedge[7] = (in[7] == 0) && (in[7] != 0);

// VERILOG-EVAL: endmodule not found
