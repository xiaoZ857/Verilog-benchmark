
module TopModule (
  input wire a,
  input wire b,
  output wire out
);

  // NOR logic: out = ~ (a | b)
  assign out = ~(a | b);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
