
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
reg currState; // Declare variable 'currState'
assign out;    // Declare output 'out' outside always block

always @(posedge clk or posedge reset) begin
    if (reset) begin
        currState <= B; // Reset the state to B when reset is active-high
        out <= 1;      // Output is 1 during reset
    end else begin
        case (currState)
            B: begin
                if (in == 0) begin
                    currState <= A;
                    out <= 1;
                end else if (in == 1) begin
                    currState <= B;
                    out <= 1;
                end
            end
            A: begin
                if (in == 0) begin
                    currState <= B;
                    out <= 0;
                end else if (in == 1) begin
                    currState <= A;
                    out <= 0;
                end
            end
        endcase
    end
end

endmodule
