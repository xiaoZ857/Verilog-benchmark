

module TopModule (
  input clk,
  input load,
  input [511:0] data,
  output reg [511:0] q
);



// VERILOG-EVAL: endmodule not found
