
module TopModule (
  input clk,
  input reset,
  output shift_ena
);
always @(posedge clk) begin
  if (reset)
    shift_ena <= 1'b1; // Reset: assert shift_ena for 4 cycles
  else if (counter == 4'b0001) // If counter is at its initial value, increment it
    counter <= counter + 1'b1;
  else if (counter > 4'b0001) // If counter is greater than its initial value, decrement it
    counter <= counter - 1'b1;
end

always @(posedge clk) begin
  if (!reset && counter < 4'b0001) // If we are not in reset and the counter is less than 4, assert shift_ena as 0
    shift_ena <= 1'b0;
end

// timescale directive should be outside of any module definition
`timescale 1ns / 1ps

reg counter = 4'b0001; // Initialize counter to 1000 (4 in binary)

// Your module interface is already provided, so I didn't include it here.

endmodule
