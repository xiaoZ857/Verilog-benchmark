
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);
logic [3:0] state;
logic [3:0] next_state;

assign start_shifting = (state == 4'b1011);

always @(posedge clk or posedge reset) begin
    if (reset)
        state <= 4'd0;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        4'd0: if (data) next_state = 4'd1; else next_state = 4'd0;
        4'd1: if (data) next_state = 4'd3; else next_state = 4'd2;
        4'd2: if (data) next_state = 4'd1; else next_state = 4'd0;
        4'd3: if (data) next_state = 4'd3; else next_state = 4'b1011;
        4'b1011: next_state = data ? 4'd3 : 4'b0010;
        default: next_state = 4'd0;
    endcase
end

endmodule
