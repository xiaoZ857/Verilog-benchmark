
module TopModule (
  input [7:0] in,
  output reg [2:0] pos
);

  always @(*) begin
    // Default to zero if no bits are high
    pos = 3'b000;
    
    // Check each bit from LSB to MSB
    if (in[0]) begin
      pos = 3'b000; // Bit position 0
    end else if (in[1]) begin
      pos = 3'b001; // Bit position 1
    end else if (in[2]) begin
      pos = 3'b010; // Bit position 2
    end else if (in[3]) begin
      pos = 3'b011; // Bit position 3
    end else if (in[4]) begin
      pos = 3'b100; // Bit position 4
    end else if (in[5]) begin
      pos = 3'b101; // Bit position 5
    end else if (in[6]) begin
      pos = 3'b110; // Bit position 6
    end else if (in[7]) begin
      pos = 3'b111; // Bit position 7
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
