

module TopModule (
  input [15:0] scancode,
  output reg left,
  output reg down,
  output reg right,
  output reg up
);



// VERILOG-EVAL: endmodule not found
