
module TopModule (
  input clk,
  input reset,
  output [3:1] ena,
  output reg [15:0] q
);
    reg [3:0] digit0, digit1, digit2, digit3;
    
    always @(posedge clk) begin
        if (reset) begin
            digit0 <= 4'b0;
            digit1 <= 4'b0;
            digit2 <= 4'b0;
            digit3 <= 4'b0;
        end
        else begin
            // Ones digit increments every clock
            if (digit0 == 4'd9) begin
                digit0 <= 4'b0;
            end
            else begin
                digit0 <= digit0 + 4'b1;
            end
            
            // Tens digit increments when ones digit wraps
            if (ena[1]) begin
                if (digit1 == 4'd9) begin
                    digit1 <= 4'b0;
                end
                else begin
                    digit1 <= digit1 + 4'b1;
                end
            end
            
            // Hundreds digit increments when tens digit wraps
            if (ena[2]) begin
                if (digit2 == 4'd9) begin
                    digit2 <= 4'b0;
                end
                else begin
                    digit2 <= digit2 + 4'b1;
                end
            end
            
            // Thousands digit increments when hundreds digit wraps
            if (ena[3]) begin
                if (digit3 == 4'd9) begin
                    digit3 <= 4'b0;
                end
                else begin
                    digit3 <= digit3 + 4'b1;
                end
            end
        end
    end
    
    // Generate enable signals
    assign ena[1] = (digit0 == 4'd9);
    assign ena[2] = (digit1 == 4'd9) && ena[1];
    assign ena[3] = (digit2 == 4'd9) && ena[2];
    
    // Combine digits into output
    always @(*) begin
        q = {digit3, digit2, digit1, digit0};
    end
endmodule
