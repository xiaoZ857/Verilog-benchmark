
// Concatenate and Split Input Vectors to Output Vectors

module TopModule (
    input [4:0] a,
    input [4:0] b,
    input [4:0] c,
    input [4:0] d,
    input [4:0] e,
    input [4:0] f,
    
    output reg [7:0] w,
    output reg [7:0] x,
    output reg [7:0] y,
    output reg [7:0] z
);

// Shift input vectors 24 bits to the left for vector concatenation
assign w = ({a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1});
reg [28:0] temp;
temp = {{a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1}};
assign w = {temp[24:20], temp[19:15]};

assign x = {{a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1}};
reg [28:0] temp_x;
temp_x = {{a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1}};
assign x = {temp_x[24:20], temp_x[19:15], temp_x[14:10], temp_x[9:5]};

reg [28:0] temp_y;
temp_y = {{a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1}};
assign y = {temp_y[24:20], temp_y[19:15], temp_y[14:10]};

reg [28:0] temp_z;
temp_z = {{a[4], b[4], c[4], d[4], e[4], f[4], 1'b1, 1'b1}};
assign z = {temp_z[24:20], temp_z[19:15]};

endmodule

// VERILOG-EVAL: errant inclusion of module definition
