
module TopModule (
    input wire clk,
    input wire [7:0] d,
    input wire reset,
    output reg [7:0] q
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        // Synchronous reset to zero
        q <= 8'b00000000;
    end else begin
        // On positive edge of clock, load the input data
        q <= d;
    end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
