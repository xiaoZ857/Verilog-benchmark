
module TopModule (
  input [99:0] in,
  output reg [99:0] out
);

always @* begin
  // Reverse the bit order
  out[99] = in[0];
  out[98] = in[1];
  out[97] = in[2];
  out[96] = in[3];
  out[95] = in[4];
  out[94] = in[5];
  out[93] = in[6];
  out[92] = in[7];
  out[91] = in[8];
  out[90] = in[9];
  out[89] = in[10];
  out[88] = in[11];
  out[87] = in[12];
  out[86] = in[13];
  out[85] = in[14];
  out[84] = in[15];
  out[83] = in[16];
  out[82] = in[17];
  out[81] = in[18];
  out[80] = in[19];
  out[79] = in[20];
  out[78] = in[21];
  out[77] = in[22];
  out[76] = in[23];
  out[75] = in[24];
  out[74] = in[25];
  out[73] = in[26];
  out[72] = in[27];
  out[71] = in[28];
  out[70] = in[29];
  out[69] = in[30];
  out[68] = in[31];
  out[67] = in[32];
  out[66] = in[33];
  out[65] = in[34];
  out[64] = in[35];
  out[63] = in[36];
  out[62] = in[37];
  out[61] = in[38];
  out[60] = in[39];
  out[59] = in[40];
  out[58] = in[41];
  out[57] = in[42];
  out[56] = in[43];
  out[55] = in[44];
  out[54] = in[45];
  out[53] = in[46];
  out[52] = in[47];
  out[51] = in[48];
  out[50] = in[49];
  out[49] = in[50];
  out[48] = in[51];
  out[47] = in[52];
  out[46] = in[53];
  out[45] = in[5

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
