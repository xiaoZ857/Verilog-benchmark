
module TopModule (
  input a,
  input b,
  output out
);

  // Implementing the AND gate logic
  assign out = a & b;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
