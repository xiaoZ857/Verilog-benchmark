
module TopModule (
  input clk,
  input reset,
  input [3:1] s,
  output reg fr3,
  output reg fr2,
  output reg fr1,
  output reg dfr
);
always @(posedge clk) begin
  if (reset) begin
    fr3 <= 1'b1;
    fr2 <= 1'b1;
    fr1 <= 1'b1;
    dfr <= 1'b1;
  end else begin
    if (s[1] == 1'b0 && s[2] == 1'b0 && s[3] == 1'b0) begin
      fr3 <= 1'b1;
      fr2 <= 1'b1;
      fr1 <= 1'b1;
      dfr <= 1'b1;
    end else if (s[1] == 1'b0 && s[2] == 1'b0 && s[3] == 1'b1) begin
      fr3 <= 1'b0;
      fr2 <= 1'b1;
      fr1 <= 1'b0;
      dfr <= 1'b0;
    end else if (s[1] == 1'b0 && s[2] == 1'b1 && s[3] == 1'b0) begin
      fr3 <= 1'b0;
      fr2 <= 1'b0;
      fr1 <= 1'b1;
      dfr <= 1'b0;
    end else if (s[1] == 1'b1 && s[2] == 1'b0 && s[3] == 1'b0) begin
      fr3 <= 1'b0;
      fr2 <= 1'b0;
      fr1 <= 1'b0;
      dfr <= 1'b1;
    end else if (s[1] == 1'b0 && s[2] == 1'b1 && s[3] == 1'b1) begin
      fr3 <= 1'b0;
      fr2 <= 1'b0;
      fr1 <= 1'b1;
      dfr <= 1'b1;
    end else if (s[1] == 1'b1 && s[2] == 1'b1 && s[3] == 1'b1) begin
      fr3 <= 1'b0;
      fr2 <= 1'b1;
      fr1 <= 1'b1;
      dfr <= 1'b1;
    end
  end
endmodule
