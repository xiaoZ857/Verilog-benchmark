
module TopModule (
  output zero
);


// VERILOG-EVAL: endmodule not found
