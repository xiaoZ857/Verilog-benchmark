

module TopModule (
  input mode,
  input too_cold,
  input too_hot,
  input fan_on,
  output heater,
  output aircon,
  output fan
);

always @(posedge clk) begin
    if (mode == 1'b1) begin // Heating mode
        heater <= too_cold;
        aircon <= 1'b0;
    end else begin // Cooling mode
        heater <= 1'b0;
        aircon <= too_hot;
    end

    fan <= (heater | aircon | fan_on);
endmodule
