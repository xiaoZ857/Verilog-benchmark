
module TopModule (
  input a,
  input b,
  output out_assign,
  output reg out_alwaysblock
);


// VERILOG-EVAL: endmodule not found
