
module TopModule (
  input clk,
  input x,
  input [2:0] y,
  output reg Y0,
  output reg z
);
reg [2:0] next_state_x0 [5]; // Changed array size to 5
reg [2:0] next_state_x1 [3];

always @(posedge clk) begin
  if (x) begin
    Y0 <= y;
    next_state_x1 <= {3'b0, 3'b0, 3'b0}; // Initialize to all zeros for first clock cycle
  end
  else begin
    Y0 <= next_state_x0[(int)y]; // Assign next state based on current state and x=0
    next_state_x1 <= {3'b0, 3'b0, 3'b0}; // Reset next_state_x1 for the next clock cycle
  end
end

always @(posedge clk) begin
  if (!x) begin
    next_state_x0 <= {3'b0, 3'b0, 3'b0, 3'b0, 3'b0}; // Initialize to all zeros for first clock cycle
  end
  else begin
    case (y)
      3'b000: next_state_x0[0] = 3'b000;
      3'b001: next_state_x0[1] = 3'b001;
      3'b010: next_state_x0[2] = 3'b010;
      3'b011: next_state_x0[3] = 3'b001;
      3'b100: next_state_x0[4] = 3'b011;
      default: next_state_x0[5] = 3'b000; // Default state for invalid input y
    endcase
  end
end

always @(posedge clk) begin
  z <= (y == 3'b100)? 1'b1 : 1'b0; // Output function for z based on current state
end

// `timescale directive should be placed outside the module definition.
`timescale 1ns / 1ps

endmodule
