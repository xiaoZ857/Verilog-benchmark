
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output q
);
assign q = (c & ~d) | (b & ~a) | (c & b);
endmodule
