

module TopModule (
  input clk,
  input d,
  output reg q
);



// VERILOG-EVAL: endmodule not found
