
module TopModule (
  input a,
  input b,
  output out_and,
  output out_or,
  output out_xor,
  output out_nand,
  output out_nor,
  output out_xnor,
  output out_anotb
);

  // Assign each output to the corresponding logic gate operation

  assign out_and = a & b;       // AND gate: a and b
  assign out_or = a | b;        // OR gate: a or b
  assign out_xor = a ^ b;       // XOR gate: a xor b
  assign out_nand = ~(a & b);   // NAND gate: a nand b
  assign out_nor = ~(a | b);    // NOR gate: a nor b
  assign out_xnor = ~(a ^ b);   // XNOR gate: a xnor b
  assign out_anotb = a & ~b;    // AND-NOT gate: a and-not b

endmodule

// VERILOG-EVAL: errant inclusion of module definition
