
module TopModule (
  input clk,
  input areset,
  input predict_valid,
  input predict_taken,
  output logic [31:0] predict_history,

  input train_mispredicted,
  input train_taken,
  input [31:0] train_history
);

reg [31:0] predict_history_reg;
reg [31:0] train_history_reg;

always @(posedge clk) begin
  if (areset) begin
    predict_history_reg <= 32'd0;
    train_history_reg <= 32'd0;
  end else if (predict_valid && !predict_taken) begin
    predict_history_reg <= predict_history_reg[31:1];
  end else if (train_mispredicted) begin
    predict_history_reg <= train_history_reg;
  end else if (train_taken) begin
    predict_history_reg <= {predict_history_reg[31:2], train_taken};
  end else begin
    predict_history_reg <= predict_history_reg[31:1];
  end

  if (train_mispredicted && !train_taken) begin
    train_history_reg <= train_history_reg[31:1] | train_taken;
  end else if (train_taken) begin
    train_history_reg <= {train_history_reg[31:2], train_taken};
  end else begin
    train_history_reg <= train_history_reg[31:1];
  end
end

assign predict_history = predict_history_reg;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
