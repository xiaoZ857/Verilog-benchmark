
module TopModule (
  input [5:0] y,
  input w,
  output Y1,
  output Y3
);

  // Logic for Y1
  assign Y1 = y[5] & w;

  // Logic for Y3
  assign Y3 = (y[4] & ~w) | (y[3] & ~w) | (y[2] & ~w) | (y[0] & ~w);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
