
module TopModule (
  input wire a,
  input wire b,
  input wire c,
  input wire d,
  input wire e,
  output [24:0] out
);

assign out[0] = ~e & e; // out[0] = e^e

wire temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14, temp15, temp16, temp17, temp18, temp19, temp20, temp21, temp22, temp23;

assign temp1 = ~a & a; // temp1 = a^a
assign temp2 = ~b & b; // temp2 = b^b
assign temp3 = ~c & c; // temp3 = c^c
assign temp4 = ~d & d; // temp4 = d^d
assign temp5 = ~e & e; // temp5 = e^e

assign out[1] = temp1; // out[1] = a^a
assign out[2] = temp2; // out[2] = b^b
assign out[3] = temp3; // out[3] = c^c
assign out[4] = temp4; // out[4] = d^d
assign out[5] = temp5; // out[5] = e^e

assign temp6 = ~a & b; // temp6 = a^b
assign temp7 = ~b & c; // temp7 = b^c
assign temp8 = ~c & d; // temp8 = c^d
assign temp9 = ~d & e; // temp9 = d^e

assign out[6] = temp6; // out[6] = a^b
assign out[7] = temp7; // out[7] = b^c
assign out[8] = temp8; // out[8] = c^d
assign out[9] = temp9; // out[9] = d^e

assign temp10 = ~a & c; // temp10 = a^c
assign temp11 = ~b & d; // temp11 = b^d
assign temp12 = ~c & e; // temp12 = c^e

assign out[10] = temp10; // out[10] = a^c
assign out[11] = temp11; // out[11] = b^d
assign out[12] = temp12; // out[12] = c^e

assign temp13 = ~a & d; // temp13 = a^d
assign temp14 = ~b & e; // temp14 = b^e

assign out[13] = temp13; // out[13] = a^d
assign out[14] = temp14; // out[14] = b^e

assign temp15 = ~c & d; // temp15 = c^d
assign temp16 = ~d & e; // temp16 = d^e

assign out[15] = temp15; // out[15] = c^d
assign out[16] = temp16; // out[16] = d^e

assign temp17 = ~a & b; // temp17 = a^b
assign temp18 = ~b & c; // temp18 = b^c
assign temp19 = ~c & d; // temp19 = c^d
assign temp20 = ~d & e; // temp20 = d^e

assign out[17] = temp17; // out[17] = a^b
assign out[18] = temp18; // out[18] = b^c
assign out[19] = temp19; // out[19] = c^d
assign out[20] = temp20; // out[20] = d^e

assign temp21 = ~a & c; // temp21 = a^c
assign temp22 = ~b & d; // temp22 = b^d
assign temp23 = ~c & e; // temp23 = c^e

assign out[2

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
