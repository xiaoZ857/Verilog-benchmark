
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);
always @(*) begin
  case (y)
    3'b000: Y2 = 0;  // State A: next state is B(001) or A(000), both have y[2]=0
    3'b001: Y2 = 1;  // State B: next state is C(010) or D(011), both have y[2]=1
    3'b010: Y2 = w;  // State C: on 0→E(100), on 1→D(011), so y[2]=w
    3'b011: Y2 = 0;  // State D: next state is F(101) or A(000), both have y[2]=0
    3'b100: Y2 = w;  // State E: on 0→E(100), on 1→D(011), so y[2]=w
    3'b101: Y2 = 1;  // State F: next state is C(010) or D(011), both have y[2]=1
    default: Y2 = 1'bx;
  endcase
end

endmodule
