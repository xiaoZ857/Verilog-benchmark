
module TopModule (
  input a,
  input b,
  input sel,
  output out
);


// VERILOG-EVAL: endmodule not found
