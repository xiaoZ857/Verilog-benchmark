

module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);



// VERILOG-EVAL: endmodule not found
