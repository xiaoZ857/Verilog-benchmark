
module TopModule (
  input clk,
  input d,
  input r,
  output logic q
);

  always_ff @(posedge clk) begin
    if (r) begin
      q <= 1'b0; // Synchronous reset to 0
    end else begin
      q <= d; // Capture the data on rising edge of clock
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
