

module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);

module FullAdder (
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

assign sum = a ^ b ^ cin;
assign cout = (a & b) | (cin & sum);

endmodule

module TopModule (
  input [3:0] x,
  input [3:0] y,
  output reg [4:0] sum,
  output reg overflow
);

wire [3:0] cin;
FullAdder fa0 (x[0], y[0], cin[0], sum[0], overflow);
FullAdder fa1 (x[1], y[1], cin[0], sum[1], cin[1]);
FullAdder fa2 (x[2], y[2], cin[1], sum[2], cin[2]);
FullAdder fa3 (x[3], y[3], cin[2], sum[3], cin[3]);

always @(posedge clk)
  overflow <= cin[3];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
