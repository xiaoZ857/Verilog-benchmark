

module TopModule (
  output one
);

assign one = 1;
endmodule
