
module TopModule (
  input [2:0] in,
  output [1:0] out
);
assign out[1] = in[2];
assign out[0] = in[1] & ~in[2];

// VERILOG-EVAL: endmodule not found
