
      ab
 cd   01  00  10  11
 00 | d | 0 | 1 | 1 |
 01 | 0 | 0 | d | d |
 11 | 0 | 1 | 1 | 1 |
 10 | 0 | 1 | 1 | 1 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
