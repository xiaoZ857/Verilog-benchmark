
module TopModule (
  input clk,
  input L,
  input q_in,
  input r_in,
  output reg Q
);


// VERILOG-EVAL: endmodule not found
