
module TopModule (
  input [2:0] in,
  output [1:0] out
);
always @(posedge clk) begin
    reg [1:0] out_reg;
    case (in)
        3'b000: out_reg <= 2'b00; // 0 ones
        3'b001: out_reg <= 2'b01; // 1 one
        3'b010: out_reg <= 2'b01; // 1 one
        3'b011: out_reg <= 2'b10; // 2 ones
        3'b100: out_reg <= 2'b01; // 1 one
        3'b101: out_reg <= 2'b10; // 2 ones
        3'b110: out_reg <= 2'b10; // 2 ones
        default: out_reg <= 2'b11; // 3 ones (for 3'b111)
    endcase
    assign out = out_reg;
end

// VERILOG-EVAL: endmodule not found
