
// Define the module that controls the cellphone's ring and vibration motors
module TopModule(
    // Inputs
    input ring,  // Indicates an incoming call
    input vibrate_mode,  // Indicates if the phone is in vibrate mode

    // Outputs
    output ringer,  // Signal to turn on the ringer
    output motor    // Signal to turn on the vibration motor
) {
    // Use the positive edge of the clock signal (clk)
    always @(posedge clk) begin
        // If an incoming call is detected and the phone is not in vibrate mode:
        if(ring && !vibrate_mode) begin
            ringer <= 1;     // Turn on the ringer
            motor <= 0;      // Turn off the vibration motor
        end else if (!ring && vibrate_mode) begin
            ringer <= 0;     // Turn off the ringer
            motor <= 1;      // Turn on the vibration motor
        end else if (ring && vibrate_mode) begin
            ringer <= 0;     // Turn off the ringer
            motor <= 1;      // Turn on the vibration motor
        end else if (!ring && !vibrate_mode) begin
            ringer <= 0;     // Turn off the ringer
            motor <= 0;      // Turn off the vibration motor
        end
    end

    // Default value for outputs
    assign default: ringer = 1'b0;
    assign default: motor = 1'b0;
}

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
