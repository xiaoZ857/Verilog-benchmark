
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output reg out
);

always @(*) begin

// VERILOG-EVAL: endmodule not found
