
module TopModule (
  input in1,
  input in2,
  output logic out
);
assign out = a & b; endmodule

// VERILOG-EVAL: endmodule not found
