
module TopModule (
  output out
);


// VERILOG-EVAL: endmodule not found
