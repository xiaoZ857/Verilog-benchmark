
module TopModule (
  input clk,
  input areset,
  input predict_valid,
  input predict_taken,
  output logic [31:0] predict_history,

  input train_mispredicted,
  input train_taken,
  input [31:0] train_history
);

  // Internal register to hold the branch history
  always_ff @(posedge clk or posedge areset) begin
    if (areset) begin
      // Asynchronous reset to zero
      predict_history <= 32'b0;
    end else if (train_mispredicted) begin
      // Load new history on misprediction
      predict_history <= {train_history, train_taken};
    end else if (predict_valid) begin
      // Shift in `predict_taken` when a valid prediction is made
      predict_history <= {predict_history[30:0], predict_taken};
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
