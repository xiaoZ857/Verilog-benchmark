
//=====================================================================
//  TopModule
//
//  Description:
//      Splits a 16‑bit input half‑word into two 8‑bit bytes.
//
//      out_hi  <= in[15:8]   // upper byte
//      out_lo  <= in[7:0]    // lower byte
//
//  Notes:
//      • The circuit is combinational – no clock or reset signals are
//        used.
//      • All signals are treated as positive‑edge triggered (i.e.
//        they update immediately on a change of 'in').
//
//=====================================================================

module TopModule (
    input  wire [15:0] in,      // 16‑bit half‑word input
    output wire [7:0]  out_hi,  // upper byte (bits 15‑8)
    output wire [7:0]  out_lo   // lower byte (bits 7‑0)
);

    // Directly map the requested slices of the input
    assign out_hi = in[15:8];
    assign out_lo = in[7:0];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
