
module TopModule (
  input clk,
  input reset,
  input s,
  input w,
  output reg z
);

reg [1:0] state;
reg [1:0] cycle_count;
reg [1:0] ones_count;
parameter A = 2'b00, B = 2'b01;

always @(posedge clk) begin
  if (reset) begin
    state <= A;
    z <= 1'b0;
    cycle_count <= 2'b00;
    ones_count <= 2'b00;
  end
  else begin
    case (state)
      A: begin
        if (s) begin
          state <= B;
          cycle_count <= 2'b00;
          ones_count <= w;
          z <= 1'b0;
        end
        else begin
          state <= A;
          z <= 1'b0;
        end
      end
      
      B: begin
        if (cycle_count == 2'b10) begin
          z <= (ones_count == 2'b10) ? 1'b1 : 1'b0;
          cycle_count <= 2'b00;
          ones_count <= w;
        end
        else begin
          cycle_count <= cycle_count + 1;
          ones_count <= ones_count + w;
          z <= 1'b0;
        end
      end
      
      default: begin
        state <= A;
        z <= 1'b0;
      end
    endcase
  end
end

endmodule
