
                x[2]x[1]
    x[4]x[3]   00   01   11   10
        00 | d | 0 | d | d |
        01 | 0 | d | 1 | 0 |
        11 | 1 | 1 | d | d |
        10 | 1 | 1 | 0 | d |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
