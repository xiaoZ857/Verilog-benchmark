
module TopModule (
  input clk,
  input in,
  input reset,
  output done
);
  // States
  localparam IDLE = 2'b00;
  localparam START = 2'b01;
  localparam DATA = 2'b10;
  localparam STOP = 2'b11;
  
  reg [1:0] state, next_state;
  reg [3:0] bit_cnt;        // Count 0-7 for 8 data bits
  reg [7:0] shift_reg;      // Shift in data bits LSB first
  reg done_reg;
  
  // State register
  always @(posedge clk) begin
    if (reset) begin
      state <= IDLE;
      bit_cnt <= 4'b0;
      shift_reg <= 8'b0;
      done_reg <= 1'b0;
    end else begin
      state <= next_state;
      
      // Bit counter and shift register updates
      case (next_state)
        IDLE: begin
          bit_cnt <= 4'b0;
          shift_reg <= 8'b0;
          done_reg <= 1'b0;
        end
        START: begin
          bit_cnt <= 4'b0;
          done_reg <= 1'b0;
        end
        DATA: begin
          // Shift in current 'in' as LSB
          shift_reg <= {in, shift_reg[7:1]};
          bit_cnt <= bit_cnt + 1;
          done_reg <= 1'b0;
        end
        STOP: begin
          // If stop bit is correct (in == 1), we can set done for one cycle
          done_reg <= (in == 1'b1);
        end
        default: begin
          bit_cnt <= bit_cnt;
          shift_reg <= shift_reg;
          done_reg <= 1'b0;
        end
      endcase
    end
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      IDLE: begin
        if (in == 1'b0)          // Start bit detected (active low)
          next_state = START;
        else
          next_state = IDLE;
      end
      START: begin
        // Wait one cycle after start bit, then go to DATA
        next_state = DATA;
      end
      DATA: begin
        if (bit_cnt == 4'd8)     // After 8 bits received
          next_state = STOP;
        else
          next_state = DATA;
      end
      STOP: begin
        if (in == 1'b1)          // Good stop bit
          next_state = IDLE;
        else                     // Missing stop bit, wait here until in==1
          next_state = STOP;
      end
      default: next_state = IDLE;
    endcase
  end
  
  assign done = done_reg;
endmodule
