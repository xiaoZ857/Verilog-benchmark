
module TopModule (
  input clk,
  input resetn,
  input x,
  input y,
  output f,
  output g
);

reg [2:0] state, next_state;
reg f_reg, g_reg;

// State encoding
parameter A = 3'b000;
parameter B = 3'b001;
parameter C = 3'b010;
parameter D = 3'b011;
parameter E = 3'b100;
parameter F = 3'b101;
parameter G = 3'b110;
parameter H = 3'b111;

// State register
always @(posedge clk) begin
  if (!resetn) begin
    state <= A;
    f_reg <= 0;
    g_reg <= 0;
  end else begin
    state <= next_state;
    case (state)
      A: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      B: begin
        f_reg <= 1;
        g_reg <= 0;
      end
      C: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      D: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      E: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      F: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      G: begin
        f_reg <= 0;
        g_reg <= 1;
      end
      H: begin
        f_reg <= 0;
        g_reg <= 0;
      end
      default: begin
        f_reg <= 0;
        g_reg <= 0;
      end
    endcase
  end
end

// Next state logic
always @(*) begin
  next_state = state;
  case (state)
    A: next_state = B;
    B: next_state = C;
    C: next_state = (x == 1) ? D : C;
    D: next_state = (x == 0) ? E : D;
    E: next_state = (x == 1) ? F : C;
    F: next_state = (y == 1) ? G : H;
    G: next_state = G;  // Stay in G permanently (g = 1)
    H: next_state = H;  // Stay in H permanently (g = 0)
    default: next_state = A;
  endcase
end

// Output assignments
assign f = f_reg;
assign g = g_reg;

endmodule
