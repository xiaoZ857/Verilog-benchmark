
module TopModule (
  input [15:0] scancode,
  output reg left,
  output reg down,
  output reg right,
  output reg up
);
always @(*) begin
    left = (scancode == 16'hE06B);
    down = (scancode == 16'hE072);
    right = (scancode == 16'hE074);
    up = (scancode == 16'hE075);
end
endmodule
