
      x[1]x[2]
      00   01   11   10
x[3]x[4]
00 |  1    0    0    1 |
01 |  0    0    0    0 |
11 |  1    1    1    0 |
10 |  1    1    0    1 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
