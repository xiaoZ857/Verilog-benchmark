

module TopModule (
  input clk,
  input resetn,
  input [1:0] byteena,
  input [15:0] d,
  output reg [15:0] q
);

always @(posedge clk or negedge resetn) begin
  if (!resetn) begin
    q <= 0;
  end else begin
    q <= d;
  end
end

always @(posedge clk) begin
  if (byteena[1]) begin
    q[15:8] <= d[15:8];
  end
  if (byteena[0]) begin
    q[7:0] <= d[7:0];
  end
end

endmodule
