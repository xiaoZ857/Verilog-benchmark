
// TopModule.v
`timescale 1ns / 1ps

module TopModule (
    input  [2:0] a,
    input  [2:0] b,
    output [2:0] out_or_bitwise,
    output       out_or_logical,
    output [5:0] out_not
);

    // Bit‑wise OR of the two 3‑bit vectors
    assign out_or_bitwise = a | b;

    // Logical OR of the two vectors (true if any bit of a or b is 1)
    assign out_or_logical = |a | |b;   // equivalent to  |(a | b)

    // Inverse of b in the upper half, inverse of a in the lower half
    assign out_not = {~b, ~a};

endmodule

// VERILOG-EVAL: errant inclusion of module definition
