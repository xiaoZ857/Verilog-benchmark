
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out_sop,
  output out_pos
);

// Sum-of-Products (SOP) for the logic-1 conditions: 2, 7, and 15
out_sop <= ~(a & b & ~c & ~d) | // 0010 (4)
         ~(a & b & c & ~d) |    // 0110 (6)
         ~(a & b & c & d) |    // 0111 (7)
         a & ~b & c & d;       // 1001 (9)

// Product-of-Sum (POS) for the logic-0 conditions: 0, 1, 4, 5, 6, 9, 10, 13, and 14
out_pos <= a & b & c & d |    // 0001 (1)
         ~a & b & c & d |     // 1001 (9)
         a & ~b & c & d |     // 1011 (13)
         a & b & ~c & d |     // 0101 (5)
         a & b & c & ~d |     // 0111 (7)
         a & b & ~c & ~d;     // 0011 (3)

// Exclude the input conditions for numbers 3, 8, 11, and 12
out_pos <= out_pos & ~(a^b^c^d);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
