
module TopModule (
  input clk,
  input areset,

  input predict_valid,
  input [6:0] predict_pc,
  output predict_taken,
  output [6:0] predict_history,

  input train_valid,
  input train_taken,
  input train_mispredicted,
  input [6:0] train_history,
  input [6:0] train_pc
);
module gshare_branch_predictor (
    input clk, // Positive clock edge
    input asreset, // Asynchronous reset active-high

    input predict_valid,
    input [6:0] predict_pc,
    output predict_taken,
    output [6:0] predict_history,

    input train_valid,
    input train_taken,
    input train_mispredicted,
    input [6:0] train_history,
    input [6:0] train_pc
);

    reg [7:0] global_branch_history;
    reg [7:0] pattern_history[127:0];
    reg [7:0] pc_hash;
    reg [4:0] history_index;

    // Gshare hash function (xor of 7-bit PC and hash of global branch history)
    assign pc_hash = predict_pc ^ global_branch_history;

    // Index into pattern history table
    always @(posedge clk) 
        begin
            if (!train_valid && !train_taken && train_mispredicted == 0)
                history_index <= {history_index[4:1], predict_pc[2]};

            else if (train_valid && !train_taken && train_mispredicted == 0)
                history_index <= {history_index, predict_pc};

            else if (train_valid && train_taken && train_mispredicted == 0)
                global_branch_history <= global_branch_history;

            else 
                begin
                    if (!predict_valid) // If training takes precedence, use the last write of global branch history
                        global_branch_history <= {history_index[4:1], predict_pc[2]};

                    else // Otherwise update pattern history table and recover branch history register
                        begin
                            pattern_history[pc_hash] <= global_branch_history;
                            if (train_taken) 
                                global_branch_history <= train_history;
                            else
                                global_branch_history <= {history_index[4:1], predict_pc[2]};
                        end

                    // Predict taken
                    predict_taken <= !!(pattern_history[pc_hash] == train_taken);

                    // Update prediction history register based on training precedence
                    predict_history <= global_branch_history;

                end
        end

    always @(posedge clk)
        if (!areset) 
            begin
                global_branch_history <= 0;
                pattern_history[127:0] <= 0;
                pc_hash <= 0;
                history_index <= 7'0;
            end

endmodule
