
x3 | x2 | x1 | f
--------------
0  | 0  | 0  | 0
0  | 0  | 1  | 0
0  | 1  | 0  | 1
0  | 1  | 1  | 1
1  | 0  | 0  | 0
1  | 0  | 1  | 1
1  | 1  | 0  | 0
1  | 1  | 1  | 1

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
