
module TopModule (
  input clk,
  input [7:0] d,
  input reset,
  output reg [7:0] q
);
always @(posedge clk) begin
    if (reset) begin
        q <= 8'b00110100;
    end else begin
        q <= d;
    end
end
endmodule
