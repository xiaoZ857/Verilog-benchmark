
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

reg [1:0] state; // State of the Lemming (00 = walking left, 01 = walking right)
reg [1:0] prev_state; // Previous state of the Lemming
reg [1:0] ground_prev; // Previous value of ground
reg [1:0] dig_prev; // Previous value of dig

// Initialize states and previous values on reset
always @(reset) begin
  state <= 2; // Walking left on reset
  prev_state <= 2;
  ground_prev <= 0;
  dig_prev <= 0;
end

// Update state based on current inputs
always @(posedge clk or negedge areset) begin
  if (areset) begin
    state <= 2; // Reset to walking left
    prev_state <= 2;
    ground_prev <= 0;
    dig_prev <= 0;
  end else begin
    // Update previous values
    ground_prev <= ground;
    dig_prev <= dig;

    // Update state based on current inputs
    if (ground == 1) begin
      if (dig == 1 && prev_state == 2) begin // Digging and walking left
        state <= 3; // Walking right while digging
      end else if (prev_state == 2) begin // Walking left
        state <= 2; // Continue walking left
      end else if (ground_prev == 0 && dig_prev == 1) begin // Falling and digging
        state <= 4; // Fall
      end else if (dig_prev == 1) begin // Digging
        state <= 3; // Walking right while digging
      end else if (bump_left == 1 && prev_state == 2) begin // Bumped on left while walking left
        state <= 1; // Walking right
      end else if (bump_right == 1 && prev_state == 1) begin // Bumped on right while walking right
        state <= 0; // Walking left
      end else if (ground_prev == 0 && bump_left == 1 && bump_right == 1) begin // Bumped on both sides while falling
        state <= 4; // Fall
      end else if (bump_left == 1 && ground_prev == 1) begin // Bumped on left while walking right
        state <= 0; // Walking left
      end else if (bump_right == 1 && ground_prev == 1) begin // Bumped on right while walking left
        state <= 1; // Walking right
      end else if (ground_prev == 1 && dig_prev == 1) begin // Digging and walking right
        state <= 3; // Walking right while digging
      end else if (dig_prev == 1) begin // Digging
        state <= 3; // Walking right while digging
      end else if (bump_left == 1 && ground_prev == 0) begin // Bumped on left while falling
        state <= 4; // Fall
      end else if (bump_right == 1 && ground_prev == 0) begin // Bumped on right while falling
        state <= 4; // Fall
      end else if (ground_prev == 0 && dig_prev == 0) begin // Falling and not digging
        state <= 4; // Fall
      end else if (bump_left == 1 && ground_prev == 1) begin // Bumped on left while walking right
        state <= 0; // Walking left
      end else if (bump_right == 1 && ground_prev == 1) begin // Bumped on right while walking left
        state <= 1; // Walking right
      end else if (ground_prev == 1 && dig_prev == 0) begin // Digging and walking right
        state <= 3; // Walking right while digging
      end else if (dig_prev == 0) begin // Not digging
        state <= 2; // Walking left
      end
    end else if (ground == 0) begin // Falling
      if (dig == 1 && prev_state == 3) begin // Digging and walking right while digging
        state <= 4; // Fall
      end else if (prev_state == 3) begin // Walking right while digging
        state <= 3; // Continue walking right while digging
      end else if (dig == 1 && prev_state == 2) begin // Digging and walking

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
