
          a
   bc | 0 | 1 |
   ----|---|---|
   00  | 0 | 1 |
   01  | 1 | 1 |
   11  | 1 | 1 |
   10  | 1 | 1 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
