

module TopModule (
  input [255:0] in,
  input [7:0] sel,
  output  out
);



// VERILOG-EVAL: endmodule not found
