
module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);

wire [1:0] nextState; // Next state of the state machine

always @(posedge clk or reset) begin
    if (reset == 1) begin      // Reset active-high, resets to OFF state
        nextState <= 2'b00;
    else if ((j == 1 && k == 0) || (k == 1)) begin
        nextState <= 2'b10;       // Transition from OFF or ON state to OFF state
    else if (j == 0) begin        // Transition within the OFF state
        nextState <= 2'b00;
    else if (j == 1 && k == 1) begin
        nextState <= 2'b01;       // Transition within the ON state
    end
end

assign out = nextState[0];   // Output is the next state in binary format

endmodule

// VERILOG-EVAL: errant inclusion of module definition
