
module TopModule (
  input clk,
  input enable,
  input S,
  input A,
  input B,
  input C,
  output reg Z
);
  reg [7:0] Q;

  always @(posedge clk) begin
    if (enable) begin
      Q[7:1] <= Q[7:2];
      Q[0] <= S;
    end
  end

  always @(*) begin
    case (A * 8 + B * 2 + C)
      0: Z = Q[0];
      1: Z = Q[1];
      2: Z = Q[2];
      3: Z = Q[3];
      4: Z = Q[4];
      5: Z = Q[5];
      6: Z = Q[6];
      7: Z = Q[7];
      default: Z = 0; // Default case to avoid latching
    endcase
  end

endmodule
