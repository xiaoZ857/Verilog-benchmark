
module TopModule (
  input clk,
  input slowena,
  input reset,
  output reg [3:0] q
);
always @(posedge clk) begin
    if (reset)
        q <= 4'b0000;
    else if (slowena)
        case (q)
            4'd9: q <= 4'b0000;
            default: q <= q + 1'b1;
        endcase
end
endmodule
