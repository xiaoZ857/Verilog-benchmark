
module TopModule (
  input clk,
  input reset,
  input data,
  output reg shift_ena,
  output reg counting,
  input done_counting,
  output reg done,
  input ack
);
always @(posedge clk) begin
    if (reset) begin
        shift_ena <= 1'b0;
        counting <= 1'b0;
        done <= 1'b0;
        state <= S_IDLE;
        pattern_reg <= 4'b0;
        shift_count <= 2'b0;
    end else begin
        case (state)
            S_IDLE: begin
                shift_ena <= 1'b0;
                counting <= 1'b0;
                done <= 1'b0;
                pattern_reg <= {pattern_reg[2:0], data};
                if (pattern_reg == 4'b1101) begin
                    state <= S_SHIFT;
                    shift_count <= 2'b0;
                    shift_ena <= 1'b1;
                end
            end
            S_SHIFT: begin
                shift_count <= shift_count + 1;
                if (shift_count == 2'b11) begin
                    shift_ena <= 1'b0;
                    counting <= 1'b1;
                    state <= S_COUNT;
                end
            end
            S_COUNT: begin
                if (done_counting) begin
                    counting <= 1'b0;
                    done <= 1'b1;
                    state <= S_DONE;
                end
            end
            S_DONE: begin
                if (ack) begin
                    done <= 1'b0;
                    state <= S_IDLE;
                    pattern_reg <= 4'b0;
                end
            end
            default: state <= S_IDLE;
        endcase
    end
end

reg [1:0] state;
reg [1:0] shift_count;
reg [3:0] pattern_reg;

localparam S_IDLE = 2'b00,
           S_SHIFT = 2'b01,
           S_COUNT = 2'b10,
           S_DONE = 2'b11;

endmodule
