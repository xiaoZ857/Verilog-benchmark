
module TopModule (
  input a,
  input b,
  output q
);


// VERILOG-EVAL: endmodule not found
