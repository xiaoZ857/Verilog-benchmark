
// Module to always output a LOW signal
module TopModule (
  // Output port for the LOW signal
  output logic zero
);

  // No inputs needed in this case, always LOW output
endmodule

// VERILOG-EVAL: errant inclusion of module definition
