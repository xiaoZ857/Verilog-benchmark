
module TopModule (
  input [99:0] in,
  output reg [98:0] out_both,
  output reg [99:1] out_any,
  output reg [99:0] out_different
);

reg [2:0] left_bit_left, right_bit_left, left_bit_right;

always_comb begin
  // Initialize signal variables based on input and their neighbours
  if (in[98] == in[99])
    left_bit_left = {1'b1, '0', '0'};
  else
    left_bit_left = {1'b0, '0', '0'};

  if (in[2] == in[1])
    right_bit_right = {1'b1, '0', '0'};
  else
    right_bit_right = {1'b0, '0', '0'};

  if (in[0] == in[99])
    left_bit_right = {1'b0, '0', '1'};
  else
    left_bit_right = {1'b1, '1', '0'};

end

assign out_both = left_bit_left;
assign out_any = right_bit_right;

always_comb begin
  // Set output signal based on difference between adjacent bits
  if (in[98] == in[99])
    out_different[98:2] = {1'b0, left_bit_left[1], left_bit_left[2]};
  else if (left_bit_left[1] == '1')
      out_different[98:2] = {1'b1, left_bit_left[1], left_bit_left[2]};
  else
    out_different[98:2] = left_bit_left;

end

always_comb begin
  // Set output signal based on difference between adjacent bits
  if (in[0] == in[99])
      out_different[100:97] = {out_different[100], right_bit_right[1], right_bit_right[2]};
  else if (right_bit_right[1] == '1')
    out_different[100:97] = {out_different[100], right_bit_right[1], right_bit_right[2]};
  else
    out_different[100:97] = right_bit_right;

end

always_comb begin
    // Set output signal based on difference between adjacent bits
      if (in[98] == in[99])
        out_different[99] = left_bit_left[0];
      else if (left_bit_left[0] == '1')
            out_different[99] = left_bit_left[0];
      else
        out_different[99] = left_bit_left[0];

end

assign out_any[100:98] = out_different[100:98];

endmodule;

// VERILOG-EVAL: errant inclusion of module definition
