
module TopModule (
  input clk,
  input areset,
  input load,
  input ena,
  input [3:0] data,
  output reg [3:0] q
);

  always @(posedge clk or posedge areset) begin
    if (areset) begin
      // Asynchronous reset to zero
      q <= 4'b0000;
    end else begin
      if (load) begin
        // Load the shift register with data
        q <= data;
      end else if (ena) begin
        // Shift right operation, shifting out from q[0]
        q <= {1'b0, q[3:1]};
      end
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
