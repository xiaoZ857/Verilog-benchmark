
module TopModule (
  input [4:0] a,
  input [4:0] b,
  input [4:0] c,
  input [4:0] d,
  input [4:0] e,
  input [4:0] f,
  output [7:0] w,
  output [7:0] x,
  output [7:0] y,
  output [7:0] z
);
  assign w = a;
  assign x = b;
  assign y = c;
  assign z = {d, e, f, 2'b11};

// VERILOG-EVAL: endmodule not found
