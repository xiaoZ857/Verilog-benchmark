
module TopModule (
  output out
);
assign out = !all_inputs;

// VERILOG-EVAL: endmodule not found
