
module TopModule (
  input [2:0] in,
  output [1:0] out
);
The Verilog module TopModule calculates

// VERILOG-EVAL: endmodule not found
