
module TopModule(
    output out
);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
