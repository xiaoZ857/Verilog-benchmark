
module TopModule (
  input clk,
  input a,
  output reg q
);
always @(posedge clk) begin
    if (a == 0) begin
        q <= 1;
    end else if (a == 1) begin
        q <= ~q; // Toggle q
    end
end

endmodule
