

module TopModule (
  input clk,
  input reset,
  input w,
  output z
);



// VERILOG-EVAL: endmodule not found
