
// This sets the simulation time scale to nanoseconds
`timescale 1ns / 1ps

module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);

always @(posedge clk) begin
  if (reset == 1) begin
    q <= 0;
  end else begin
    if (q == 9) begin
      q <= 0;
    end else begin
      q <= q + 1;
    end
  end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
