
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out_sop,
  output out_pos
);

// Minimum Sum-of-Products (SOP) form for out_sop
assign out_sop = (~a & ~b & ~c & ~d) | 
                 (~a & ~b & c & d) | 
                 (~a & b & ~c & d) |
                 (~a & b & c & ~d) |
                 (a & ~b & ~c & d) |
                 (a & ~b & c & ~d) |
                 (a & b & ~c & ~d);

// Minimum Product-of-Sums (POS) form for out_pos
assign out_pos = (~a | ~b | ~c | ~d) &
                (~a | ~b | c | d) &
                (~a | b | ~c | d) &
                (~a | b | c | ~d) &
                (a | ~b | ~c | d) &
                (a | ~b | c | ~d) &
                (a | b | ~c | ~d);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
