
module TopModule (
  input x,
  input y,
  output z
);
assign z = x == 1'b0 && y == 1'b0;
endmodule
