
module TopModule (
  input a,
  input b,
  output sum,
  output cout
);


// VERILOG-EVAL: endmodule not found
