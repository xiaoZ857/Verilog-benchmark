
// Shift the input vector to the right by one position and select the last bit
assign o0 = vec[2];

// Select the least significant bit of the input vector
assign o1 = vec[1];

// Select the middle bit of the input vector
assign o2 = vec[0];

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
