
module TopModule (
  input wire a,
  input wire b,
  input wire c,
  input wire d,
  output wire q
);

assign q = (!a && !b && !c && !d) || ((!a && !b && !c && d) && ((!a && b) || (a && c))) || ((!a && b && c && !d) && ((!b && c) || (b && d)));

endmodule

// VERILOG-EVAL: errant inclusion of module definition
