
module TopModule (
    input clk,
    input [7:0] in,
    input reset,
    output done
);

    reg [2:0] state;
    reg [7:0] message_in;
    wire [7:0] out;

    reg [3:0] done_state; // New variable to track the state of the done signal

    always @(posedge clk) begin
        if (reset) begin
            state <= 3'b000; // Reset to idle state
            message_in <= 8'b0; // Clear message buffer
            done_state <= 4'b0000; // Reset done state
        end else begin
            message_in <= in[2:0]; // Update message buffer with new byte

            case(state)
                3'b000: // Idle state
                    if (message_in[3] == 1) begin
                        state <= 3'b001; // Start of message detected
                        done_state <= 4'b0000; // Reset done state
                    end
                3'b001: // Message start detected, waiting for second byte
                    if (message_in[2] == 1) begin
                        state <= 3'b010; // Second byte received, waiting for third byte
                        done_state <= 4'b0000; // Reset done state
                    end else begin
                        state <= 3'b000; // Invalid message, reset to idle state
                        done_state <= 4'b0000; // Reset done state
                    end
                3'b010: // Message in progress, waiting for third byte
                    if (message_in[1] == 1) begin
                        state <= 3'b011; // Third byte received, signal done
                        done_state <= 4'b1111; // Signal done
                    end else begin
                        state <= 3'b000; // Invalid message, reset to idle state
                        done_state <= 4'b0000; // Reset done state
                    end
                default: // Invalid state
                    state <= 3'b000;
            endcase

            if (done_state == 4'b1111) begin // Done state
                done <= 1'b1;
                state <= 3'b000; // Reset to idle state after done signal is sent
                done_state <= 4'b0000; // Reset done state
            else begin
                done <= 1'b0;
            end
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
