
module TopModule (
  input [5:0] y,
  input w,
  output reg Y1,
  output reg Y3
);

assign Y1 = y[1]; // Y1 is the input of state flip-flop y[1]
assign Y3 = (y[3] || (w && (~y[0] & ~y[2]))); // Y3 is the input of state flip-flop y[3]

always @(posedge clk) begin
  if (Y1) begin
    case ({Y1, Y3})
      2'b00: Y1 <= 0;
      2'b01: Y1 <= 1;
      2'b10: Y1 <= 0; // A state

      2'b11: if (Y3) begin
                Y3 <= 0;
              end else begin
                Y3 <= 1;
              end; // B state
    end

    case ({Y1, ~Y3})
      2'b00: Y1 <= 0;
      2'b01: Y1 <= 0;
      2'b10: Y1 <= 0; // A state

      2'b11: if (w) begin
                Y3 <= 0;
              end else begin
                Y3 <= 1;
              end; // D state

    case ({Y3})
      2'b0: begin
        if (Y3) begin
          case ({Y1})
            2'b0: Y1 <= 1; // C state
            2'b1: Y1 <= 0; // D state
          end
        end else begin
          case ({Y1})
            2'b0: Y1 <= 0; // A state
            2'b1: Y1 <= 1; // B state
          end
        end
    end

    case ({~Y3})
      2'b0: begin
        if (w) begin
          case ({Y1})
            2'b0: Y1 <= 1; // E state
            2'b1: Y1 <= 0; // D state
          end
        end else begin
          case ({Y1})
            2'b0: Y1 <= 0; // A state
            2'b1: Y1 <= 1; // B state
          end
        end
    end

    case ({Y1, ~w})
      2'b00: Y1 <= 1; // F state
      2'b01: Y1 <= 0; // D state
    endcase
  end
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
