
module TopModule (
  input clk,
  input load,
  input [511:0] data,
  output reg [511:0] q
);
always @(posedge clk) begin
    if (load)
        q <= data;
    else begin
        q[0] <= 1'b0; // Boundary condition, always off
        q[511] <= 1'b0; // Boundary condition, always off
        for (int i = 1; i < 511; i++) begin
            q[i] <= q[i-1] ^ q[i+1];
        end
    end
end
endmodule
