
module TopModule (
  input clk,
  input j,
  input k,
  input reset,
  output out
);
  // Define the states
  parameter OFF = 2'b00;
  parameter ON  = 2'b01;

  // Declare the state register
  reg current_state;
  reg out;

  // Assign the output based on the current state
  always @(current_state) begin
    case (current_state)
      OFF: out = 0;
      ON : out = 1;
      default: out = 0;  // Default case for safety
    endcase
  end

  // Synchronous reset
  always @(posedge clk) begin
    if (reset) begin
      current_state <= OFF;
    end else begin
      // State transition logic
      case (current_state)
        OFF: begin
          if (j) begin
            current_state <= ON;
          end else begin
            current_state <= OFF;
          end
        end
        ON: begin
          if (k) begin
            current_state <= OFF;
          end else begin
            current_state <= ON;
          end
        end
        default: current_state <= OFF; // Safety net
      endcase
    end
  end

endmodule
