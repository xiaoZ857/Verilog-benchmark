
module TopModule (
  input clock,
  input a,
  output reg p,
  output reg q
);
always @(posedge clock) begin
    // Update p with the current value of a at each clock cycle
    p <= a;
    
    // Check if a was 1 in the last cycle to update q accordingly
    if (last_a == 1'b1) begin
        q <= p; // Capture the current value of p when last_a was 1
    end else begin
        q <= 1'b0; // Reset q to 0 otherwise
    end
    
    // Store the current value of a for use in the next cycle
    last_a <= a;
end

// Additional register needed to store the previous state of 'a'
reg last_a;

initial begin
    last_a = 1'b0; // Initialize last_a at the start
end

endmodule
