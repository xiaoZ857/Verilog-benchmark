
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
