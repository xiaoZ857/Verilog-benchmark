

module TopModule (
  input clk,
  input reset,
  input in,
  output disc,
  output flag,
  output err
);



// VERILOG-EVAL: endmodule not found
