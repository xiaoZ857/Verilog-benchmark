
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);


// VERILOG-EVAL: endmodule not found
