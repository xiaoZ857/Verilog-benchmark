

module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  output walk_left,
  output walk_right
);

 ```verilog
always @(posedge clk or negedge areset)
begin
    if (areset)
        walk_left <= 1'b1;
        walk_right <= 1'b0;
    else if (bump_left && !walk_left)
        walk_left <= 1'b0;
        walk_right <= 1'b1;
    else if (bump_right && !walk_right)
        walk_left <= 1'b0;
        walk_right <= 1'b1;
    else
        walk_left <= walk_left;
        walk_right <= !walk_left;
end

assign walk_left = walk_left ^ walk_right; // Ensure only one output is high at any given time

endmodule

// VERILOG-EVAL: abnormal backticks count
