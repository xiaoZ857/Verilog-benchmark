

module TopModule (
  input clk,
  input reset,
  output shift_ena
);

reg [3:0] state; // FSM state variables
always @(posedge clk or posedge reset) begin
  if (reset) begin
    state <= 4'b0001; // Reset state, assert shift_ena for 4 cycles
  end else begin
    case (state)
      4'b0001: state <= 4'b0010; // Move to next state
      4'b0010: state <= 4'b0100; // Move to next state
      4'b0100: state <= 4'b1000; // Move to next state
      4'b1000: state <= 4'b0001; // Reset back to initial state, shift_ena is always asserted during this state
    default: state <= 4'b0000; // Invalid state, reset FSM
    endcase
  end
end

assign shift_ena = (state == 4'b0001) || (state == 4'b0010) || (state == 4'b0100) || (state == 4'b0100); // shift_ena is asserted during the first 4 states

endmodule
