
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);
reg [2:0] state, next_state;

localparam
    IDLE_LEFT     = 3'b000,
    WALK_RIGHT    = 3'b001,
    WALK_LEFT     = 3'b010,
    FALL          = 3'b011,
    DIG           = 3'b100;

assign aaah = (state == FALL);
assign digging = (state == DIG);

always @(posedge areset or posedge clk) begin
    if (areset)
        state <= IDLE_LEFT;
    else
        state <= next_state;
end

always @(*) begin
    case (state)
        IDLE_LEFT: begin
            if (~ground)
                next_state = FALL;
            else if (bump_left)
                next_state = WALK_RIGHT;
            else if (dig && ground)
                next_state = DIG;
            else
                next_state = IDLE_LEFT;
        end

        WALK_RIGHT: begin
            if (~ground)
                next_state = FALL;
            else if (bump_right || bump_left)
                next_state = WALK_LEFT;
            else if (dig && ground)
                next_state = DIG;
            else
                next_state = WALK_RIGHT;
        end

        WALK_LEFT: begin
            if (~ground)
                next_state = FALL;
            else if (bump_right || bump_left)
                next_state = WALK_RIGHT;
            else if (dig && ground)
                next_state = DIG;
            else
                next_state = WALK_LEFT;
        end

        FALL: begin
            if (ground)
                next_state = state == IDLE_LEFT ? IDLE_LEFT :
                             state == WALK_RIGHT ? WALK_RIGHT :
                             WALK_LEFT;
            else
                next_state = FALL;
        end

        DIG: begin
            if (~ground)
                next_state = FALL;
            else
                next_state = DIG;
        end

        default: next_state = IDLE_LEFT;
    endcase
end

always @(*) begin
    case (state)
        IDLE_LEFT: begin
            walk_left = 1'b1;
            walk_right = 1'b0;
        end
        
        WALK_RIGHT: begin
            walk_left = 1'b0;
            walk_right = 1'b1;
        end

        WALK_LEFT: begin
            walk_left = 1'b1;
            walk_right = 1'b0;
        end

        FALL, DIG: begin
            walk_left = (state == IDLE_LEFT || state == WALK_LEFT);
            walk_right = (state == IDLE_LEFT) ? 1'b0 : (state == WALK_RIGHT) ? 1'b1 : 1'b0;
        end
        
        default: begin
            walk_left = 1'b0;
            walk_right = 1'b0;
        end
    endcase
end

endmodule
