
module TopModule (
  input [31:0] in,
  output [31:0] out
);
  // Internal signals to hold the reversed bytes
  wire [7:0] byte0;
  wire [7:0] byte1;
  wire [7:0] byte2;
  wire [7:0] byte3;

  // Extract individual bytes from the input
  assign byte0 = in[7:0];
  assign byte1 = in[15:8];
  assign byte2 = in[23:16];
  assign byte3 = in[31:24];

  // Construct the output with reversed byte order
  assign out = {byte3, byte2, byte1, byte0};

endmodule
