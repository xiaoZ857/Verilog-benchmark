
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out,
  output out_n
);
  wire and1_out;
  wire and2_out;

  // First layer: Two AND gates
  and1_out = a & b;
  and2_out = c & d;

  // Second layer: OR gate and NOT gate
  out = and1_out | and2_out;
  out_n = ~out;

endmodule
