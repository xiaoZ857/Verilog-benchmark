
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
  // Define states
  parameter A = 2'b00
  parameter B = 2'b01

  // State register
  reg current_state;

  // Output register
  reg out;

  // Synchronous reset
  always @(posedge clk or posedge areset) begin
    if (areset) begin
      current_state <= B;
    end else begin
      case (current_state)
        A: begin
          if (in == 0) begin
            current_state <= B;
          end else begin
            current_state <= A;
          end
        end
        B: begin
          if (in == 0) begin
            current_state <= B;
          end else begin
            current_state <= B;
          end
        end
        default: begin
          current_state <= B; // Default to B in case of unexpected state
        end
      endcase
    end
  end

  // Output logic (Moore machine)
  always @(current_state) begin
    case (current_state)
      A: out = 1;
      B: out = 0;
      default: out = 0; // Default output
    endcase
  end

endmodule
