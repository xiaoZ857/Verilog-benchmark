
module TopModule (
  input in,
  output out
);

  // Directly assign the input to the output
  assign out = in;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
