
module TopModule (
  output zero
);
  zero = 1'b0;
endmodule
