
module TopModule (
  input clk,
  input [7:0] d,
  input reset,
  output reg [7:0] q
);

  // Declare an array of D flip-flops
  reg [7:0] dff_q;

  // Synchronous reset logic
  always @(posedge clk) begin
    if (reset) begin
      q <= 0;
    end else begin
      q <= d;
    end
  end

endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
