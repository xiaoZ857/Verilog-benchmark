
module TopModule (
  input clk,
  input reset,
  input x,
  output reg z
);
always @(posedge clk) begin
  if (reset) begin
    z <= 1'b0;
  end else begin
    case (y[2:0])
      3'b000: begin
        if (x == 1'b0)
          y <= 3'b000;
        else
          y <= 3'b001;
      end
      3'b001: begin
        if (x == 1'b0)
          y <= 3'b001;
        else
          y <= 3'b100;
      end
      3'b010: begin
        if (x == 1'b0)
          y <= 3'b010;
        else
          y <= 3'b001;
      end
      3'b011: begin
        if (x == 1'b0)
          y <= 3'b001;
        else
          y <= 3'b010;
        z <= 1'b1;
      end
      3'b100: begin
        if (x == 1'b0)
          y <= 3'b011;
        else
          y <= 3'b100;
        z <= 1'b1;
      end
      default: begin
        y <= 3'b000;
      end
    endcase
  end
end

endmodule
