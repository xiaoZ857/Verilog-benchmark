
module TopModule (
  input [4:1] x,
  output logic f
);
always @(*) begin
  if ((x[1] == 1'b0 && x[2] == 1'b0) && (x[3] == 1'b0 && x[4] == 1'b0))
    f = 1'b0;
  else if ((x[1] == 1'b0 && x[2] == 1'b1) && (x[3] == 1'b0 && x[4] == 1'b1))
    f = 1'b0;
  else if ((x[1] == 1'b1 && x[2] == 1'b1 && x[3] == 1'b1 && x[4] == 1'b1))
    f = 1'b1;
  else if ((x[1] == 1'b1 && x[2] == 1'b1 && x[3] == 1'b1 && x[4] == 1'b0))
    f = 1'b1;
  else
    f = 1'b0;
endmodule
