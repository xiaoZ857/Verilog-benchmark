
// TopModule.v
// 3‑bit pass‑through + split into 3 single‑bit outputs
module TopModule (
    input  wire [2:0] vec,  // 3‑bit input vector
    output wire [2:0] outv, // same vector as output
    output wire       o2,   // vec[2]
    output wire       o1,   // vec[1]
    output wire       o0    // vec[0]
);

// Combinational assignments – no clock needed
assign outv = vec;      // forward the whole vector
assign o0   = vec[0];   // split out bit 0
assign o1   = vec[1];   // split out bit 1
assign o2   = vec[2];   // split out bit 2

endmodule

// VERILOG-EVAL: errant inclusion of module definition
