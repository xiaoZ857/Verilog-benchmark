

module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);

  reg [1:0] current_state;
  reg [1:0] next_state;

  always @(posedge clk or negedge aresetn) begin
    if (!aresetn) begin
      current_state <= 0;
      z <= 0;
    end else begin
      current_state <= next_state;
    end
  end

  always @(*) begin
    next_state = current_state;
    case (current_state)
      2'b00: begin
        if (x) begin
          next_state = 2'b01;
        end else begin
          next_state = 2'b00;
        end
      end
      2'b01: begin
        if (!x) begin
          next_state = 2'b00;
        end else begin
          next_state = 2'b01;
        end
      end
      2'b10: begin
        if (x) begin
          next_state = 2'b01;
        end else begin
          next_state = 2'b10;
        end
      end
      default: begin
        next_state = 2'b00;
      end
    endcase

    if (current_state == 2'b10 && x) begin
      z = 1;
    end else begin
      z = 0;
    end
  end
endmodule
