
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
