
module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);

  always @(posedge clk) begin
    if (reset) begin
      q <= 32'h1;
    end else begin
      // Galois LFSR with taps at positions 32, 22, 2, and 1
      // Feedback bit is the LSB (q[0])
      q[31] <= q[30] ^ q[0];  // Position 32 tap
      q[30] <= q[29];
      q[29] <= q[28];
      q[28] <= q[27];
      q[27] <= q[26];
      q[26] <= q[25];
      q[25] <= q[24];
      q[24] <= q[23];
      q[23] <= q[22] ^ q[0];  // Position 22 tap
      q[22] <= q[21];
      q[21] <= q[20];
      q[20] <= q[19];
      q[19] <= q[18];
      q[18] <= q[17];
      q[17] <= q[16];
      q[16] <= q[15];
      q[15] <= q[14];
      q[14] <= q[13];
      q[13] <= q[12];
      q[12] <= q[11];
      q[11

// VERILOG-EVAL: endmodule not found
