

module TopModule (
  input in,
  input [9:0] state,
  output [9:0] next_state,
  output out1,
  output out2
);



// VERILOG-EVAL: endmodule not found
