
module TopModule (
  output zero
);

  assign zero = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
