

module TopModule (
  input x,
  input y,
  output z
);



// VERILOG-EVAL: endmodule not found
