
module TopModule (
  input p1a,
  input p1b,
  input p1c,
  input p1d,
  input p1e,
  input p1f,
  output p1y,
  input p2a,
  input p2b,
  input p2c,
  input p2d,
  output p2y
);

  wire and1_out;
  wire and2_out;

  // p1y is the OR of two 3-input AND gates
  assign and1_out = p1a & p1b & p1c;
  assign and2_out = p1d & p1e & p1f;
  assign p1y = and1_out | and2_out;

  // p2y is the OR of two 2-input AND gates
  assign p2y = (p2a & p2b) | (p2c & p2d);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
