
// ------------------------------------------------------------
//  TopModule
//  ---------
//  Implements a 2‑input AND gate in two different ways:
//
//      1)  Continuous assignment (wire)
//      2)  Combinational always block (reg)
//
//  The module has no clock – all logic is purely combinational.
// ------------------------------------------------------------
`timescale 1ns/1ps

module TopModule (
    input  wire a,                // first AND input
    input  wire b,                // second AND input
    output wire out_assign,       // result from continuous assignment
    output reg  out_alwaysblock   // result from always block
);

// ------------------------------------------------------------
// 1) Continuous assignment
// ------------------------------------------------------------
assign out_assign = a & b;

// ------------------------------------------------------------
// 2) Combinational always block
// ------------------------------------------------------------
always @(*) begin
    out_alwaysblock = a & b;
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
