
module TopModule (
  output out
);
// Assign 0 to the output 'out' at the beginning of simulation
initial begin
  out = 0;
end

// VERILOG-EVAL: endmodule not found
