
module TopModule (
  input a,
  input b,
  output out_assign,
  output reg out_alwaysblock
);

  // Continuous assignment using assign statement
  assign out_assign = a & b;

  // Combinational logic using always block
  always @(*) begin
    out_alwaysblock = a & b;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
