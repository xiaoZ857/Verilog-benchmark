

module TopModule (
  input clk,
  input reset,
  input [31:0] in,
  output reg [31:0] out
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        out <= 32'b0; // Reset the output to zero
    end else begin
        for (int i = 0; i < 32; i++) begin
            if ((in[i] == 1'b1) && (~in[i + 1] == 1'b0)) begin
                out[i] <= 1'b1; // Set the output to 1 for the transition bit
            end
        end
    end
end

always @(posedge clk) begin
    out <= out; // Propagate the values in the output register
end

assign out_sync = reset | (~reset & out); // Provide a synchronous output for use elsewhere

endmodule
