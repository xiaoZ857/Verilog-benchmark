
module TopModule (
  input clk,
  input a,
  input b,
  output q,
  output state
);
logic state_reg;

always @(posedge clk) begin
  state_reg <= state_reg;
end

always @(posedge clk) begin
  if (a == 1 && b == 1 && state_reg == 0) begin
    state_reg <= 1;
  end else if (a == 0 && b == 0 && state_reg == 1) begin
    state_reg <= 0;
  end else if (a == 1 && b == 0 && state_reg == 1) begin
    state_reg <= 0;
  end else if (a == 0 && b == 1 && state_reg == 0) begin
    state_reg <= 1;
  end else if (a == 1 && b == 1 && state_reg == 1) begin
    state_reg <= 1;
  end else if (a == 0 && b == 0 && state_reg == 0) begin
    state_reg <= 0;
  end else if (a == 1 && b == 0 && state_reg == 0) begin
    state_reg <= 0;
  end else if (a == 0 && b == 1 && state_reg == 1) begin
    state_reg <= 0;
  end else if (a == 1 && b == 0 && state_reg == 1) begin
    state_reg <= 0;
  end
end

assign q = state_reg;
assign state = state_reg;
endmodule
