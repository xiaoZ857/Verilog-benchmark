
module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);
always @(posedge clk) begin
  if (reset) begin
    q <= 5'b11111;  // Reset to all 1s
  end else begin
    // Galois LFSR shifting right
    q[4] <= q[3] ^ q[0];  // Bit 5 (position 5) has tap
    q[3] <= q[4];         // Bit 4 shifts right
    q[2] <= q[1] ^ q[0];  // Bit 3 (position 3) has tap
    q[1] <= q[2];         // Bit 2 shifts right
    q[0] <= q[1];         // Bit 1 shifts right
  end
end

endmodule
