
module TopModule (
  input clk,
  input j,
  input k,
  input areset,
  output out
);


// VERILOG-EVAL: endmodule not found
