

module TopModule (
  input clk,
  input in,
  input reset,
  output done
);

  reg [2:0] state;
  reg [2:0] next_state;
  reg [2:0] bit_count;
  reg data_valid;
  reg stop_bit_expected;

  always @(posedge clk) begin
    if (reset) begin
      state <= 3'b000; // Idle state
      data_valid <= 1'b0;
      stop_bit_expected <= 1'b0;
      bit_count <= 3'b000;
      done <= 1'b0;
    end else begin
      state <= next_state;
      done <= 1'b0;
      if (state == 3'b000) begin // Idle
        if (in == 1'b0) begin
          next_state <= 3'b001; // Start bit detected
        end else begin
          next_state <= 3'b000;
        end
      end else if (state == 3'b001) begin // Start bit
        if (bit_count == 3'b000) begin
          next_state <= 3'b010; // Data bits
          bit_count <= 3'b000;
        end else begin
          next_state <= 3'b010;
        end
      end else if (state == 3'b010) begin // Data bits
        if (bit_count == 3'b111) begin // 8 data bits received
          next_state <= 3'b011; // Stop bit expected
          stop_bit_expected <= 1'b1;
        end else begin
          bit_count <= bit_count + 3'b001;
          next_state <= 3'b010;
        end
      end else if (state == 3'b011) begin // Stop bit expected
        if (in == stop_bit_expected) begin
          next_state <= 3'b000; // Back to idle
          data_valid <= 1'b1;
          done <= 1'b1;
        end else begin
          next_state <= 3'b011; // Wait for stop bit
        end
      end
    end
  end

endmodule
