
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out,
  output out_n
);


// VERILOG-EVAL: endmodule not found
