
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);
always @(posedge clk) begin
    if (reset) begin
        done <= 1'b0;
        out_byte <= 8'b0;
        state <= IDLE;
        bit_count <= 3'b0;
        shift_reg <= 8'b0;
    end else begin
        case (state)
            IDLE: begin
                done <= 1'b0;
                if (in == 1'b0) begin
                    state <= START;
                end
            end
            START: begin
                if (in == 1'b1) begin
                    state <= IDLE;
                end else begin
                    state <= DATA;
                    bit_count <= 3'b0;
                end
            end
            DATA: begin
                shift_reg <= {in, shift_reg[7:1]};
                if (bit_count == 3'b111) begin
                    state <= STOP;
                end else begin
                    bit_count <= bit_count + 1;
                end
            end
            STOP: begin
                if (in == 1'b1) begin
                    done <= 1'b1;
                    out_byte <= shift_reg;
                    state <= IDLE;
                end else begin
                    state <= START;
                end
            end
            default: state <= IDLE;
        endcase
    end
end

localparam IDLE = 2'b00;
localparam START = 2'b01;
localparam DATA = 2'b10;
localparam STOP = 2'b11;

reg [1:0] state;
reg [2:0] bit_count;
reg [7:0] shift_reg;
endmodule
