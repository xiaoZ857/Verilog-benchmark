
module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);

// Macro to calculate the neighbour cell index
#define NEIGHBOUR(i, j) ((i + 1) % 16 * 16 + (j + 1) % 16)

always @(posedge clk) begin
  if (load) begin
    q <= data;
  end else begin
    logic [255:0] new_state;

    // Iterate through all cells
    for (int i = 0; i < 16; i++) begin
      for (int j = 0; j < 16; j++) begin
        int count = 0;

        // Count the number of living neighbors
        count += q[NEIGHBOUR(i-1, j-1)] +    // top left
                 q[NEIGHBOUR(i-1, j )] +     // top center
                 q[NEIGHBOUR(i-1, j+1)] +    // top right
                 q[NEIGHBOUR( i   , j-1)] +   // current cell left
                 q[NEIGHBOUR( i   , j+1)] +   // current cell right
                 q[NEIGHBOUR(i+1, j-1)] +    // bottom left
                 q[NEIGHBOUR(i+1, j )] +     // bottom center
                 q[NEIGHBOUR(i+1, j+1)];      // bottom right

        // Update the state based on the number of neighbors
        if (count == 3 || (count == 2 && q[NEIGHBOUR(i,j)])) begin
          new_state[NEIGHBOUR(i,j)] = 1;
        end else if (count != 2) begin
          new_state[NEIGHBOUR(i,j)] = 0;
        end
      end
    end

    q <= new_state;
  end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
