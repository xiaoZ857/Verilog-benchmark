
module TopModule (
  output zero
);

  // Assign a constant LOW value to the output 'zero'
  assign zero = 1'b0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
