
    x[4] x[3] x[2] x[1] | f
    ---------------------|------
    0       0           0      1
    0       1           0      0
    1       0           1      0
    1       1           1      0
    1       1           0      1

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
