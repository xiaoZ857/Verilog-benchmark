
module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);
always @(posedge clk) begin
    if (reset) begin
        q <= 5'b00001;
    end
    else begin
        q[4] <= q[3] ^ q[0];  // Tap at position 5
        q[3] <= q[2];         // No tap, just shift
        q[2] <= q[1] ^ q[0];  // Tap at position 3
        q[1] <= q[0];         // No tap, just shift
        q[0] <= q[4];         // MSB shifts to LSB
    end
end

endmodule
