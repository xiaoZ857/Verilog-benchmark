
module TopModule (
  input in,
  input [1:0] state,
  output reg [1:0] next_state,
  output out
);
  always @(*) begin
    case (state)
      2'b00: begin // A
        if (in == 1'b0) next_state = 2'b00;
        else next_state = 2'b01;
      end
      2'b01: begin // B
        if (in == 1'b0) next_state = 2'b10;
        else next_state = 2'b01;
      end
      2'b10: begin // C
        if (in == 1'b0) next_state = 2'b00;
        else next_state = 2'b11;
      end
      2'b11: begin // D
        if (in == 1'b0) next_state = 2'b10;
        else next_state = 2'b01;
      end
      default: next_state = 2'b00;
    endcase
  end

  assign out = (state == 2'b11) ? 1'b1 : 1'b0;

endmodule
