

module TopModule (
  input clk,
  input resetn,
  input x,
  input y,
  output f,
  output g
);



// VERILOG-EVAL: endmodule not found
