

module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);

always @(posedge clk) begin
  if (reset) begin
    q <= 0;
  end else begin
    q <= q + 1;
  end
endmodule
