
module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);
// -----------------------------------------------------------------------------
//  Full‑adder helper module
// -----------------------------------------------------------------------------
module FullAdder (
    input  a,
    input  b,
    input  cin,
    output sum,
    output cout
);
    // The 2‑bit addition of a, b and cin produces a 3‑bit result.
    // The most significant bit is the carry out, the least significant bit is the sum.
    assign {cout, sum} = a + b + cin;
endmodule

// -----------------------------------------------------------------------------
//  4‑bit adder with overflow bit
// -----------------------------------------------------------------------------
    // Internal carry wires
    wire c0, c1, c2;

    // Full‑adder instantiations
    FullAdder fa0 (
        .a   (x[0]),
        .b   (y[0]),
        .cin (1'b0),
        .sum (sum[0]),
        .cout(c0)
    );

    FullAdder fa1 (
        .a   (x[1]),
        .b   (y[1]),
        .cin (c0),
        .sum (sum[1]),
        .cout(c1)
    );

    FullAdder fa2 (
        .a   (x[2]),
        .b   (y[2]),
        .cin (c1),
        .sum (sum[2]),
        .cout(c2)
    );

    FullAdder fa3 (
        .a   (x[3]),
        .b   (y[3]),
        .cin (c2),
        .sum (sum[3]),
        .cout(sum[4])   // overflow bit
    );

endmodule
