
module TopModule (
  input wire a,
  input wire b,
  output wire q
);

assign q = (a ^ b);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
