

module TopModule (
  input clk,
  input reset,
  input s,
  input w,
  output reg z
);



// VERILOG-EVAL: endmodule not found
