

module TopModule (
  input [99:0] in,
  output out_and,
  output out_or,
  output out_xor
);



// VERILOG-EVAL: endmodule not found
