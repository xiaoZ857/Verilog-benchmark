
module TopModule (
    input wire in1,
    input wire in2,
    output logic out
);

assign out = ~(in1 | in2);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
