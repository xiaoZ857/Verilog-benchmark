
module TopModule(
    input [4:1] x,
    output logic f
);

    assign f = 
        x[0] & (x[2] | ~x[3]) & (~x[1] | (x[2] & ~x[4]));

endmodule

// VERILOG-EVAL: errant inclusion of module definition
