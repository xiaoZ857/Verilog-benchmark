
module TopModule (
  input d,
  input done_counting,
  input ack,
  input [9:0] state, // 10-bit one-hot current state
  output B3_next,
  output S_next,
  output S1_next,
  output Count_next,
  output Wait_next,
  output done,
  output counting,
  output shift_ena
);
// Next-state logic
assign S_next = (state[0] & ~d) |        // S --d=0--> S
                (state[1] & ~d) |        // S1 --d=0--> S
                (state[3] & ~d) |        // S110 --d=0--> S
                (state[9] & ack);        // Wait --ack=1--> S

assign S1_next = state[0] & d;           // S --d=1--> S1

// Note: S11_next is not required as output, but needed for S110_next
// S11_next = (state[1] & d) | (state[2] & d)  // S1 --d=1--> S11, S11 --d=1--> S11

assign S110_next = state[2] & ~d;        // S11 --d=0--> S110

assign B0_next = state[3] & d;           // S110 --d=1--> B0

assign B1_next = state[4];               // B0 --always--> B1

assign B2_next = state[5];               // B1 --always--> B2

assign B3_next = state[6];               // B2 --always--> B3

assign Count_next = state[7];            // B3 --always--> Count

assign Wait_next = state[8] & done_counting; // Count --done_counting=1--> Wait

// Output logic
assign shift_ena = state[4] | state[5] | state[6] | state[7]; // B0, B1, B2, B3
assign counting = state[8]; // Count state
assign done = state[9]; // Wait state
endmodule
