
module TopModule (
    input clk,
    input reset,
    input ena,
    output reg pm,
    output reg [7:0] hh,
    output reg [7:0] mm,
    output reg [7:0] ss
);

reg [1:0] hours;
reg [3:0] tens_minutes;
reg [3:0] ones_minutes;
reg [3:0] seconds;

reg [1:0] am_pm;
reg [1:0] hour_12;
reg [1:0] minute_60;
reg [1:0] second_60;

initial begin
    // Initialize counters to 00:00:00 AM
    hours = 0;
    tens_minutes = 0;
    ones_minutes = 0;
    seconds = 0;
    
    am_pm = 0; // AM by default
    hour_12 = 1; // 12-hour clock
    minute_60 = 0; // 60-minute clock
    second_60 = 0; // 60-second clock
    
end

always @(posedge clk) begin
    if (ena && !reset) begin
        // Increment seconds, minutes, and hours on every enable pulse
        if (seconds == 59) begin
            seconds = 0;
            minute_60 = minute_60 + 1;
            if (minute_60 == 60) begin
                minute_60 = 0;
                hour_12 = hour_12 + 1;
                if (hour_12 == 13) begin // 24-hour clock
                    hour_12 = 0;
                end
            end
        end else if (minutes == 59) begin
            minutes = 0;
            second_60 = second_60 + 1;
            if (second_60 == 60) begin
                second_60 = 0;
                minute_60 = minute_60 + 1;
                if (minute_60 == 60) begin // 24-hour clock
                    minute_60 = 0;
                    hour_12 = hour_12 + 1;
                    if (hour_12 == 13) begin
                        hour_12 = 0;
                    end
                end
            end
        end else if (hours == 11) begin // 24-hour clock
            hours = 0;
            minute_60 = minute_60 + 1;
            if (minute_60 == 60) begin
                minute_60 = 0;
                hour_12 = hour_12 + 1;
                if (hour_12 == 13) begin
                    hour_12 = 0;
                end
            end
        end else begin
            hours = hours + 1;
            if (hours == 12) begin // 24-hour clock
                hours = 0;
                minute_60 = minute_60 + 1;
                if (minute_60 == 60) begin
                    minute_60 = 0;
                    hour_12 = hour_12 + 1;
                    if (hour_12 == 13) begin
                        hour_12 = 0;
                    end
                end
            end
        end
        
        // Update BCD values
        hh = hours * 16 + tens_minutes * 2 + ones_minutes;
        mm = minute_60 * 10 + second_60;
        ss = seconds;
        
    end else if (ena) begin
        // Reset counters on enable pulse when reset is active
        if (reset == 1) begin
            hours = 0;
            tens_minutes = 0;
            ones_minutes = 0;
            seconds = 0;
            
            am_pm = 0; // AM by default
            hour_12 = 1; // 12-hour clock
            minute_60 = 0; // 60-minute clock
            second_60 = 0; // 60-second clock
            
        end else begin
            // Increment seconds, minutes, and hours on every enable pulse
            if (seconds == 59) begin
                seconds = 0;
                minute_60 = minute_60 + 1;
                if (minute_60 == 60) begin
                    minute_60 = 0;
                    hour_12 = hour_12 + 1;
                    if (hour_12 == 13) begin // 24-hour clock
                        hour_12 = 0;
                    end
                end
            end else if (minutes == 59) begin
                minutes = 0;
                second_60 = second_60 + 1;
                if (second_60 == 60) begin
                    second_60 = 0;
                    minute_60 = minute_60 + 1

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
