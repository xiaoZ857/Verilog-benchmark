
module TopModule (
  input clk,
  input resetn,
  input x,
  input y,
  output f,
  output g
);
reg state = 0; // FSM state variable
wire f, g; // Declare output signals as wires since they are driven by the top module
reg last_x = 0; // Last value of x
reg last_last_x = 0; // Two clock cycles ago value of x
reg last_y = 0; // Last value of y
reg y_count = 0; // Counts the number of times y is observed to be 1 since the last reset or g transition

always @(posedge clk) begin
    if (!resetn) begin
        state <= 0; // Reset the FSM to state A
        f <= 0; // Set output f to 0 when reset
        g <= 0; // Set output g to 0 when reset
    end else begin
        case (state)
            0: begin // State A
                if (f == 0) begin
                    assign f = 1; // Assign f to 1 for one clock cycle after reset
                end
                last_last_x <= last_x; // Store the value of x from two clock cycles ago
                last_x <= x; // Store the current value of x
                if (last_x == last_last_x && last_x == 1) begin // Check if x has produced the values 1, 0, 1 in three successive clock cycles
                    state <= 1; // Transition to next state
                end
            end
            1: begin // Monitoring g and y
                last_y <= y; // Store the current value of y
                if (g == 1 && y == 1) begin // If y has the value 1, maintain g = 1 permanently
                    y_count <= 0; // Reset y_count
                end else if (g == 1 && y == 0) begin // If y does not have the value 1, set g = 0 permanently
                    assign g = 0;
                end
                if (y_count < 2 && y == 1) begin // Count the number of times y is observed to be 1 since the last reset or g transition
                    y_count <= y_count + 1;
                end
            end
        endcase
    end
end

// No need for a separate 'timescale' directive as it should already be set in your Verilog environment.

endmodule
