
module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] pedge
);
always @(posedge clk) begin
  for (int i = 0; i < 8; i++) begin
    if (!in[i] && posedge[i]) // Check for rising edge (0 to 1 transition)
      pedge[i] <= 1'b1; // Set output bit the cycle after a 0 to 1 transition occurs
  end
end

// VERILOG-EVAL: endmodule not found
