
module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);
logic [2:0] state, next_state;
assign start_shifting = (state == 3'b101);

always_ff @(posedge clk or posedge reset) begin
    if (reset)
        state <= 3'b000;
    else
        state <= next_state;
end

always_comb begin
    case (state)
        3'b000: next_state = data ? 3'b001 : 3'b000;
        3'b001: next_state = data ? 3'b010 : 3'b000;
        3'b010: next_state = data ? 3'b011 : 3'b100;
        3'b011: next_state = data ? 3'b101 : 3'b000;
        3'b100: next_state = data ? 3'b001 : 3'b000;
        3'b101: next_state = 3'b101; // Remain in this state
        default: next_state = 3'b000;
    endcase
end

endmodule
