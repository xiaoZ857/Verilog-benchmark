

module TopModule (
  input [7:0] in,
  output [7:0] out
);



// VERILOG-EVAL: endmodule not found
