
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);
 ```verilog
always @(posedge clk or posedge reset) begin
    if (reset) begin
        reg [23:0] message;
        done <= 1'b0;
    end else begin
        reg [7:0] current_byte = in;
        static int state = 0;

        always @* begin
            case (state)
                0: begin
                    if (current_byte[3]) begin
                        message <= current_byte;
                        state += 1;
                    end
                end,
                1: begin
                    message <= {message, current_byte};
                    state += 1;
                    if (state == 4) begin
                        done <= 1'b1;
                        state = 0;
                    end
                end,
                default: state = 0;
            endcase
        end

        assign out_bytes = message[23:0];
    end
end
endmodule

// VERILOG-EVAL: abnormal backticks count
