
module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);
always @(posedge clk) begin
    if (load)
        q <= data;
    else begin
        integer i, j, count;
        logic [3:0] neighbors;

        for (i = 0; i < 16; i++) begin
            for (j = 0; j < 16; j++) begin
                // Calculate the number of live neighbors
                neighbors = 0;
                
                // Check all eight possible neighbors with wrap-around using modulo operation
                neighbors += q[((i-1) + 16) % 16 * 16 + ((j-1) + 16) % 16];
                neighbors += q[((i-1) + 16) % 16 * 16 + j];
                neighbors += q[((i-1) + 16) % 16 * 16 + ((j+1) + 16) % 16];
                neighbors += q[i * 16 + ((j-1) + 16) % 16];
                neighbors += q[i * 16 + ((j+1) + 16) % 16];
                neighbors += q[((i+1) + 16) % 16 * 16 + ((j-1) + 16) % 16];
                neighbors += q[((i+1) + 16) % 16 * 16 + j];
                neighbors += q[((i+1) + 16) % 16 * 16 + ((j+1) + 16) % 16];

                // Apply the rules of the game
                if (q[i*16+j] == 0 && (neighbors == 3))
                    q[i*16+j] <= 1;
                else if (q[i*16+j] == 1 && (neighbors < 2 || neighbors > 3))
                    q[i*16+j] <= 0;
            end
        end
    end
end

endmodule
