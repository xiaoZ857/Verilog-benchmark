
//=====================================================================
//  7420 – Two 4‑input NAND gates
//
//  Module name:  TopModule
//
//  Ports
//  ├─ p1a, p1b, p1c, p1d : 4 inputs to the first NAND gate
//  │  p1y                : output of the first NAND gate
//  ├─ p2a, p2b, p2c, p2d : 4 inputs to the second NAND gate
//  │  p2y                : output of the second NAND gate
//=====================================================================
`timescale 1ns/1ps

module TopModule (
    input  wire p1a,
    input  wire p1b,
    input  wire p1c,
    input  wire p1d,
    output wire p1y,
    input  wire p2a,
    input  wire p2b,
    input  wire p2c,
    input  wire p2d,
    output wire p2y
);

    // 4‑input NAND gate #1
    assign p1y = ~(p1a & p1b & p1c & p1d);

    // 4‑input NAND gate #2
    assign p2y = ~(p2a & p2b & p2c & p2d);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
