
module TopModule (
  input clk,
  input resetn,
  input in,
  output out
);
logic [3:0] shift_reg;

always @(posedge clk) begin
  if (!resetn) begin
    shift_reg <= 0;
  end else begin
    shift_reg <= {shift_reg[3:1], in};
  end
end

assign out = shift_reg[0];

endmodule
