
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);
reg y_next [1]; // Next state of y[1] and y[0] combined in a single register

always @(posedge clk) begin
  case (y[2])
    0: y_next = w ? 3'b01 : 3'b00; // next state for A based on input w
    1: y_next = (w == 1'b0) ? 3'b00 : 3'b01; // next state for B
    2: y_next = w ? 3'b10 : 3'b01; // next state for C based on input w
    3: y_next = (w == 1'b0) ? 3'b10 : 3'b00; // next state for D
    4: y_next = w ? 3'b00 : 3'b11; // next state for E based on input w
    5: y_next = 3'b11; // next state for F is always 1
    default: y_next = 3'bx; // Unreachable state, set to 'x' (unknown) value
  endcase

  Y2 <= y[2]; // Assign current state (Y2) to output
  assign y[0] = y_next[1]; // Assign next state of y[0]
end

// VERILOG-EVAL: endmodule not found
