
module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);


// VERILOG-EVAL: endmodule not found
