
module TopModule (
  input clk,
  input reset,
  output [3:1] ena,
  output reg [15:0] q
);
always @(posedge clk) begin
  if (reset) begin
    q <= 16'h0000;
  end else begin
    // Increment ones digit always
    if (q[3:0] == 4'h9) begin
      q[3:0] <= 4'h0;
      // Enable tens digit when ones rolls over
      if (q[7:4] == 4'h9) begin
        q[7:4] <= 4'h0;
        // Enable hundreds digit when tens rolls over
        if (q[11:8] == 4'h9) begin
          q[11:8] <= 4'h0;
          // Enable thousands digit when hundreds rolls over
          if (q[15:12] == 4'h9) begin
            q[15:12] <= 4'h0;
          end else begin
            q[15:12] <= q[15:12] + 1;
          end
        end else begin
          q[11:8] <= q[11:8] + 1;
        end
      end else begin
        q[7:4] <= q[7:4] + 1;
      end
    end else begin
      q[3:0] <= q[3:0] + 1;
    end
  end
end

// Generate enable signals
assign ena[1] = (q[3:0] == 4'h9);  // Enable tens when ones is 9
assign ena[2] = (q[7:4] == 4'h9) && (q[3:0] == 4'h9);  // Enable hundreds when tens and ones are 9
assign ena[3] = (q[11:8] == 4'h9) && (q[7:4] == 4'h9) && (q[3:0] == 4'h9);  // Enable thousands when hundreds, tens, and ones are 9

endmodule
