

module TopModule (
  input a,
  input b,
  input c,
  output out
);

assign out = (a & b) | ((~a & ~b) | (~c & ~b));
endmodule
