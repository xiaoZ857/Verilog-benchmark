
module TopModule (
  input [99:0] in,
  output [98:0] out_both,
  output [99:1] out_any,
  output [99:0] out_different
);
// Continuous assignments for the required relationships
assign out_both      = in[98:0] & in[99:1];          // both current and left neighbour are 1
assign out_any       = in[99:1] | in[98:0];          // either current or right neighbour is 1
assign out_different = in ^ {in[0], in[99:1]};       // current bit differs from left neighbour (wrap‑around)
endmodule
