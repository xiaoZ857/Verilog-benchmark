
module TopModule (
  input [7:0] in,
  output reg [2:0] pos
);
Here’s a straightforward, synthesizable implementation of a **least‑significant‑bit priority encoder

// VERILOG-EVAL: endmodule not found
