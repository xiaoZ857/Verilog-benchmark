
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out,
  output out_n
);
  wire and_ab;
  wire and_cd;

  // First layer: AND gates
  and_ab = a & b;
  and_cd = c & d;

  // Second layer: OR gate and NOT gate
  or or_gate (
    .a(and_ab),
    .b(and_cd),
    .out(out)
  );

  not not_gate (
    .in(out),
    .out(out_n)
  );

endmodule
