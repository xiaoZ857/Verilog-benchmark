
assign out_and = (a & b); // AND gate
assign out_or = (a | b); // OR gate
assign out_xor = (a ^ b); // XOR gate
assign out_nand = !(a & b); // NAND gate
assign out_nor = !(a | b); // NOR gate
assign out_xnor = !(a ^ b); // XNOR gate
assign out_anotb = (a & !b); // AND-NOT gate

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
