

module TopModule (
  input clk,
  input x,
  output z
);



// VERILOG-EVAL: endmodule not found
