
module TopModule (
  input [1023:0] in,
  input [7:0] sel,
  output [3:0] out
);
assign out = (sel == 8'b00000000) ? in[3:0] :
             (sel == 8'b00000001) ? in[7:4] :
             (sel == 8'b00000010) ? in[11:8] :
             (sel == 8'b00000011) ? in[15:12] :
             (sel == 8'b00000100) ? in[19:16] :
             (sel == 8'b00000101) ? in[23:20] :
             (sel == 8'b00000110) ? in[27:24] :
             (sel == 8'b00000111) ? in[31:28] :
             (sel == 8'b00001000) ? in[35:32] :
             (sel == 8'b00001001) ? in[39:36] :
             (sel == 8'b00001010) ? in[43:40] :
             (sel == 8'b00001011) ? in[47:44] :
             (sel == 8'b00001100) ? in[51:48] :
             (sel == 8'b00001101) ? in[55:52] :
             (sel == 8'b00001110) ? in[59:56] :
             (sel == 8'b00001111) ? in[63:60] :
             (sel == 8'b00010000) ? in[67:64] :
             (sel == 8'b00010001) ? in[71:68] :
             (sel == 8'b00010010) ? in[75:72] :
             (sel == 8'b00010011) ? in[79:76] :
             (sel == 8'b00010100) ? in[83:80] :
             (sel == 8'b00010101) ? in[87:84] :
             (sel == 8'b00010110) ? in[91:88] :
             (sel == 8'b00010111) ? in[95:92] :
             (sel == 8'b00011000) ? in[99:96] :
             (sel == 8'b00011001) ? in[103:100] :
             (sel == 8'b00011010) ? in[107:104] :
             (sel == 8'b00011011) ? in[111:108] :
             (sel == 8'b00011100) ? in[115:112] :
             (sel == 8'b00011101) ? in[119:116] :
             (sel == 8'b00011110) ? in[123:120] :
             (sel == 8'b00011111) ? in[127:124] :
             (sel == 8'b00100000) ? in[131:128] :
             (sel == 8'b00100001) ? in[135:132] :
             (sel == 8'b00100010) ? in[139:136] :
             (sel == 8'b00100011) ? in[143:140] :
             (sel == 8'b00100100) ? in[147:144] :
             (sel == 8'b00100101) ? in[151:148] :
             (sel == 8'b00100110) ? in[155:152] :
             (sel == 8'b00100111) ? in[159:156] :
             (sel == 8'b00101000) ? in[163:160] :
             (sel == 8'b00101001) ? in[167:164] :
             (sel == 8'b00101010) ? in[171:168] :
             (sel == 8'b00101011) ? in[175:172] :
             (sel == 8'b00101100) ? in[179:176] :
             (sel == 8'b00101101) ? in[183:180] :
             (sel == 8'b00101110) ? in[187:184] :
             (sel == 8'b00101111) ? in[191:188] :
             (sel == 8'b00110000) ? in[195:192] :
             (sel == 8'b00110001) ? in[199:196] :
             (sel == 8'b00110010) ? in[203:200] :
             (sel == 8'b00110011) ? in[207:204] :
             (sel == 8'b00110100) ? in[211:208] :
             (sel == 8'b00110101)

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
