
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);

  // State definitions
  localparam IDLE = 2'b00;
  localparam BYTE1 = 2'b01;
  localparam BYTE2 = 2'b10;
  localparam DONE = 2'b11;
  
  // State registers
  reg [1:0] state, next_state;
  
  // Message storage registers
  reg [7:0] byte1, byte2, byte3;
  reg [23:0] out_bytes_reg;
  reg done_reg;
  
  // State transition logic
  always @(*) begin
    next_state = state;
    case (state)
      IDLE: begin
        if (in[3]) begin
          next_state = BYTE1;
        end
      end
      BYTE1: begin
        next_state = BYTE2;
      end
      BYTE2: begin
        next_state = DONE;
      end
      DONE: begin
        if (in[3]) begin
          next_state = BYTE1;
        end else begin
          next_state = IDLE;
        end
      end
    endcase
  end
  
  // Sequential logic
  always @(posedge clk) begin
    if (reset) begin
      state <= IDLE;
      byte1 <= 8'b0;
      byte2 <= 8'b0;
      byte3 <= 8'b0;
      out_bytes_reg <= 24'b0;
      done_reg <= 1'b0;
    end else begin
      state <= next_state;
      
      case (state)
        IDLE: begin
          if (in[3]) begin
            byte1 <= in;
            done_reg <= 1'b0;
          end
        end
        BYTE1: begin
          byte2 <= in;
          done_reg <= 1'b0;
        end
        BYTE2: begin
          byte3 <= in;
          out_bytes_reg <= {byte1, byte2, in};
          done_reg <= 1'b1;
        end
        DONE: begin
          if (in[3]) begin
            byte1 <= in;
            done_reg <= 1'b0;
          end else begin
            done_reg <= 1'b0;
          end
        end
      endcase
    end
  end
  
  // Output assignments
  assign out_bytes = out_bytes_reg;
  assign done = done_reg;

endmodule
