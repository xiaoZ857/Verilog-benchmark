
module TopModule (
  input clock,
  input a,
  output reg p,
  output reg q
);
always @(posedge clock) begin  
    if (a) begin 
        p <= 1'b1;  
        q <= p;
    end else begin
        q <= 1'b0;
    end
end

endmodule
