
module TopModule (
  input clk,
  input in,
  output logic out
);


// VERILOG-EVAL: endmodule not found
