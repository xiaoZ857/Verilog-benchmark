
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
  // State encoding
  localparam logic STATE_A = 1'b0;
  localparam logic STATE_B = 1'b1;

  logic state, next_state;

  // State register with asynchronous reset
  always_ff @(posedge clk or posedge areset) begin
    if (areset)
      state <= STATE_B;          // reset to state B
    else
      state <= next_state;       // normal state transition
  end

  // Next‑state logic (combinational)
  always_comb begin
    case (state)
      STATE_A: begin
        if (in == 1'b0)
          next_state = STATE_B;
        else
          next_state = STATE_A;
      end
      STATE_B: begin
        if (in == 1'b0)
          next_state = STATE_A;
        else
          next_state = STATE_B;
      end
      default: next_state = STATE_B; // safety default
    endcase
  end

  // Moore output (depends only on state)
  assign out = (state == STATE_B) ? 1'b1 : 1'b0;
endmodule
