
module TopModule (
  input [2:0] a,
  output reg [15:0] q
);


// VERILOG-EVAL: endmodule not found
