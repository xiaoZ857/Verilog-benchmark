
module TopModule (
  input clock,
  input a,
  output reg p,
  output reg q
);
reg state = 0; // 0 for State 1, 1 for State 2

always @(posedge clock) begin
  if (state === 0) begin
    if (a) begin
      q <= 1'b1;
      state <= 1'b1;
    end else begin
      p <= 1'b0;
      q <= 1'b0;
    end
  end else begin
    if (a) begin
      p <= 1'b1;
      q <= 1'b1;
    end else begin
      p <= 1'b0;
      q <= 1'b0;
      state <= 1'b0; // transition back to State 1 after a delay
    end
  end
end

// Add initial block for resetting the state to 0 at the beginning
initial begin
  #5 $finish; // Simulation ends after 5ns
  state <= 0; // Reset the state to 0 initially
end

// Timescale directive should be outside of the module definition
`timescale 1ns / 1ps

endmodule
