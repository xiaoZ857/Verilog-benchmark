
module TopModule (

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
