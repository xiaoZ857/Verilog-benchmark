
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);
  reg [23:0] out_bytes_reg;
  reg [2:0] state;
  reg done_reg;

  always @(posedge clk) begin
    if (reset) begin
      state <= 0;
      done_reg <= 0;
      out_bytes_reg <= 0;
    end else begin
      case (state)
        0: begin // Initial state - searching for first byte
          if (in[3] == 1) begin
            state <= 1;
            out_bytes_reg <= {0, in[7:0]};
          end else begin
            state <= 0;
            out_bytes_reg <= 0;
          end
        end
        1: begin // Received first byte - searching for second byte
          if (in[3] == 1) begin
            state <= 1;
            out_bytes_reg <= {0, in[7:0]};
          end else begin
            state <= 2;
            out_bytes_reg <= {{out_bytes_reg[7:0], in[7:0]}};
          end
        end
        2: begin // Received first two bytes - searching for third byte
          if (in[3] == 1) begin
            state <= 1;
            out_bytes_reg <= {0, in[7:0]};
          end else begin
            state <= 2;
            out_bytes_reg <= {{out_bytes_reg[15:0], in[7:0]}};
          end
        end
        default: begin
          state <= 0;
        end
      endcase
    end
  end

  assign out_bytes = out_bytes_reg;
  assign done = (state == 2);

// VERILOG-EVAL: endmodule not found
