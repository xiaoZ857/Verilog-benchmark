
module TopModule (
  input [1:0] A,
  input [1:0] B,
  output z
);


// VERILOG-EVAL: endmodule not found
