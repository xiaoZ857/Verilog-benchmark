
       c
     0   1
b\c | 00 | 01 |
   -------------
   0 |  0 |  1 |
a  -------------
   1 |  1 |  1 |
   -------------
   1 |  1 |  1 |

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
