

module TopModule (
  input clk,
  input shift_ena,
  input count_ena,
  input data,
  output reg [3:0] q
);



// VERILOG-EVAL: endmodule not found
