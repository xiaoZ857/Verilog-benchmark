
module TopModule (
  input clk,
  input areset,

  input predict_valid,
  input [6:0] predict_pc,
  output predict_taken,
  output [6:0] predict_history,

  input train_valid,
  input train_taken,
  input train_mispredicted,
  input [6:0] train_history,
  input [6:0] train_pc
);
reg [6:0] ghr;
reg [1:0] pht [0:127];

wire [6:0] predict_index = predict_pc ^ ghr;
wire [1:0] predict_counter = pht[predict_index];

assign predict_taken = predict_counter[1];
assign predict_history = ghr;

wire [6:0] train_index = train_pc ^ train_history;
reg [1:0] train_counter;

// PHT update logic
always @(posedge clk or posedge areset) begin
    if (areset) begin
        ghr <= 7'b0;
        // Initialize PHT to weakly not-taken (01)
        for (integer i = 0; i < 128; i = i + 1) begin
            pht[i] <= 2'b01;
        end
    end else begin
        // Training has priority over prediction updates
        if (train_valid) begin
            // Update PHT for training
            train_counter = pht[train_index];
            if (train_taken) begin
                // Saturating increment
                if (train_counter != 2'b11) begin
                    pht[train_index] <= train_counter + 1;
                end
            end else begin
                // Saturating decrement
                if (train_counter != 2'b00) begin
                    pht[train_index] <= train_counter - 1;
                end
            end

            // Recover ghr if mispredicted
            if (train_mispredicted) begin
                // ghr becomes train_history shifted with actual outcome
                ghr <= {train_history[5:0], train_taken};
            end else if (predict_valid) begin
                // Normal update with predicted direction (only if no misprediction recovery)
                ghr <= {ghr[5:0], predict_taken};
            end
        end else if (predict_valid) begin
            // Normal update with predicted direction
            ghr <= {ghr[5:0], predict_taken};
        end
    end
end
endmodule
