
module TopModule (
  input clk,
  input reset,
  output shift_ena
);
logic [3:0] counter;

always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
        counter <= 4'b1111;
        shift_ena <= 1'b1;
    end else begin
        if (counter != 4'b0000)
            counter <= counter - 1'b1;
        else
            shift_ena <= 1'b0;
    end
end

assign shift_ena = (counter != 4'b0000);

// VERILOG-EVAL: endmodule not found
