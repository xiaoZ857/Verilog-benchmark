
module TopModule (
  input [4:1] x,
  output logic f
);
assign f = (x[1:0] == 2'b00 && (x[3] ^ x[4])) || 
           (x[1:0] == 2'b11 && (x[3] | x[4] | (x[3] & x[4]))) ||
           (x[1:0] == 2'b10 && ((x[3] & ~x[4]) | (~x[3] & x[4]) | x[4])) ||
           (x[1:0] == 2'b01 && 1'b0);
endmodule
