
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out
);
assign out = (!a | b) & (!b | c) & (!c | d);

// VERILOG-EVAL: abnormal backticks count
