
module TopModule (
  input wire clk,
  input wire resetn,
  input [3:1] r,
  output reg [3:1] g
);

// State codes
parameter STATE_A = 2'b00;
parameter STATE_B = 2'b01;
parameter STATE_C = 2'b10;
parameter STATE_D = 2'b11;

// FSM state variables
reg [1:0] current_state;

always @(posedge clk or posedge resetn) begin
  if (resetn) begin
    current_state <= STATE_A;
  end else begin
    case (current_state)
      STATE_A: begin
        if (r[1] == 1) begin
          current_state <= STATE_B;
          g[1] <= 1'b1;
        end else if (r[2] == 1) begin
          current_state <= STATE_C;
          g[2] <= 1'b1;
        end else if (r[3] == 1) begin
          current_state <= STATE_D;
          g[3] <= 1'b1;
        end else begin
          current_state <= STATE_A;
        end
      end
      STATE_B: begin
        if (r[1] == 0) begin
          current_state <= STATE_A;
        end else begin
          current_state <= STATE_B;
        end
      end
      STATE_C: begin
        if (g2 && r[2] == 0) begin
          current_state <= STATE_A;
        end else begin
          current_state <= STATE_C;
        end
      end
      STATE_D: begin
        if (r[3] == 0) begin
          current_state <= STATE_A;
        end else begin
          current_state <= STATE_D;
        end
      end
    endcase
  end
end

// Continuous assignment for g[i] outputs
assign g[1] = (current_state == STATE_B);
assign g[2] = (current_state == STATE_C);
assign g[3] = (current_state == STATE_D);

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
