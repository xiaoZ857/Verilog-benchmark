
module TopModule (
  input clk,
  input resetn,
  input in,
  output out
);


// VERILOG-EVAL: endmodule not found
