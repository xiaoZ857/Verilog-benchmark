
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
always @(posedge clk or negedge areset) begin
  if (areset) begin
    // Reset the state machine to initial state B when reset is high
    A <= 1'b0;
    B <= 1'b1;
  end else begin
    assign out = B;
    case (A)
      // A transition table
      1'b0: B <= in;
      1'b1: B <= ~A;
    endcase

    case (B)
      // B transition table
      1'b0: A <= in;
      1'b1: A <= ~B;
    endcase
  end
end

reg A, B;

endmodule
