
always @ (posedge clk) begin
    case ({c, d}) // Using {c, d} as they are the most significant bits in the K-map
        2'b00: out = 1'b0; // For cd = 00
        2'b01: 
            if (c == 1'b0 && d == 1'b0) out = 1'b0;
            else out = 1'bx; // Don't care for other combinations when cd = 01
        2'b11: out = 1'b1; // For cd = 11
        2'b10: out = 1'b1; // For cd = 10
        default: out = 1'bx; // Default case for don't-care values
    endcase
end

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
