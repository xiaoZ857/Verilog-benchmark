
// 4‑state Moore machine (A,B,C,D)
// State encoding :  A = 2'b00,  B = 2'b01,  C = 2'b10,  D = 2'b11
//
//  State | Next state (in=0) | Next state (in=1) | Output
//  -------------------------------------------------------
//  A     | A                | B                | 0
//  B     | C                | B                | 0
//  C     | A                | D                | 0
//  D     | C                | B                | 1
//
//  Only the combinational logic (next_state & out) is required.

module TopModule (
    input  wire        in,          // input
    input  wire [1:0]  state,       // current state
    output reg  [1:0]  next_state,  // next state (combinational)
    output wire        out          // output
);

    // ------------------------------------------------------------
    // Output logic – Moore output depends only on the current state
    // ------------------------------------------------------------
    assign out = (state == 2'b11) ? 1'b1 : 1'b0;   // 1 only for state D

    // ------------------------------------------------------------
    // State transition logic – combinational
    // ------------------------------------------------------------
    always @(*) begin
        case (state)
            2'b00:   // State A
                next_state = in ? 2'b01 : 2'b00;   // B if in=1, else A
            2'b01:   // State B
                next_state = in ? 2'b01 : 2'b10;   // B if in=1, else C
            2'b10:   // State C
                next_state = in ? 2'b11 : 2'b00;   // D if in=1, else A
            2'b11:   // State D
                next_state = in ? 2'b01 : 2'b10;   // B if in=1, else C
            default: // safety net – stay in A
                next_state = 2'b00;
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
