
module TopModule (
  input clk,
  input d,
  output reg q
);
assign q = d; endmodule

// VERILOG-EVAL: endmodule not found
