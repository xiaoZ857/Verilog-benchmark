
module TopModule (
  input [254:0] in,
  output reg [7:0] out
);
// Count the number of '1's in the input vector
reg [7:0] count = 8'd0;
for (int i = 0; i < 255; i++) begin
    count = count + ((in[i] == 1) ? 1 : 0);
end

// Store the population count in the output signal
out = count;

endmodule
