
module TopModule (
  output zero
);
  assign zero = 1'b0;
endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
