
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);
typedef enum logic [1:0] {
    STATE_A = 2'b00,
    STATE_B = 2'b01,
    STATE_C = 2'b10,
    STATE_D = 2'b11
} state_t;

// Current and next state registers
state_t state, next_state;

// State register – synchronous with active‑high reset
always_ff @(posedge clk) begin
    if (reset)
        state <= STATE_A;          // reset to state A
    else
        state <= next_state;       // normal state transition
end

// Next‑state logic (combinational)
always_comb begin
    next_state = state;            // default: stay in current state
    case (state)
        STATE_A: next_state = (in == 1'b0) ? STATE_A : STATE_B;
        STATE_B: next_state = (in == 1'b0) ? STATE_C : STATE_B;
        STATE_C: next_state = (in == 1'b0) ? STATE_A : STATE_D;
        STATE_D: next_state = (in == 1'b0) ? STATE_C : STATE_B;
        default: next_state = STATE_A;
    endcase
end

// Output logic (Moore output)
assign out = (state == STATE_D) ? 1'b1 : 1'b0;

endmodule
