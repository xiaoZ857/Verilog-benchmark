
Y1 (next B)  = y[0] & w
Y3 (next D)  = (~w) & (y[1] | y[2] | y[4] | y[5])

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
