

module TopModule (
  output zero
);

assign zero = 0;

// VERILOG-EVAL: endmodule not found
