
module TopModule (
  input [4:1] x,
  output logic f
);
  always_comb begin
    if ((x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 1 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 1) ||
        (x[1] == 0 && x[2] == 0 && x[3] == 0 && x[4] == 0) ||
        (x[

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
