
module TopModule (
  input [7:0] in,
  output [31:0] out
);
assign out = {in[7:0], 24'd1} & {in[7:0], 24'd1};

endmodule
