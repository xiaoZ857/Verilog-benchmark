
module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);


// VERILOG-EVAL: endmodule not found
