
module TopModule (
  input in,
  input [9:0] state,
  output [9:0] next_state,
  output out1,
  output out2
);
 ```verilog
always @(posedge clk) begin
    if (in)
        case (state)
            0: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            1: begin
                next_state <= {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b1;
            end
            2: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            3: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            4: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            5: begin
                next_state <= {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            6: begin
                next_state <= {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
            7: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b1;
            end
            8: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b1;
                out2 <= 1'b0;
            end
            9: begin
                next_state <= {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                out1 <= 1'b0;
                out2 <= 1'b0;
            end
        endcase
    else
       

// VERILOG-EVAL: endmodule not found
