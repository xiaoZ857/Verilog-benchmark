
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
) {
  reg [2:0] state;
  reg [7:0] message_in;
  reg [1:0] byte_count;

  always @(posedge clk) begin
    if (reset) begin
      state <= 3'b000;
      message_in <= 8'd0;
      byte_count <= 2'b00;
    end else begin
      byte_count <= byte_count + 1;
      message_in <= in[byte_count-1:byte_count-2];

      case(state)
        3'b000: if (message_in[3] == 1) state <= 3'b001; else state <= 3'b000;
        3'b001: if (message_in[3] == 0 && byte_count == 2) done <= 1;
                  if (byte_count < 2) state <= 3'b001;
                  else state <= 3'b000;
        default: state <= 3'b000;
      endcase
    end
  end

  assign done = message_in[3] == 0 && byte_count == 2;
}
endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
