

module TopModule (
  input clk,
  input reset,
  input w,
  output z
);

  localparam STATE_A = 2'b00;
  localparam STATE_B = 2'b01;
  localparam STATE_C = 2'b10;
  localparam STATE_D = 2'b11;
  localparam STATE_E = 2'b10;
  localparam STATE_F = 2'b01;

  reg [1:0] current_state;
  reg [1:0] next_state;

  always @(posedge clk) begin
    if (reset) begin
      current_state <= STATE_A;
    else begin
      current_state <= next_state;
    end
  end

  always @(*) begin
    next_state = current_state;
    case (current_state)
      STATE_A: begin
        if (w)
          next_state = STATE_B;
        else
          next_state = STATE_A;
      end
      STATE_B: begin
        if (w)
          next_state = STATE_C;
        else
          next_state = STATE_D;
      end
      STATE_C: begin
        if (w)
          next_state = STATE_E;
        else
          next_state = STATE_D;
      end
      STATE_D: begin
        if (w)
          next_state = STATE_F;
        else
          next_state = STATE_A;
      end
      STATE_E: begin
        if (w)
          next_state = STATE_E;
        else
          next_state = STATE_D;
      end
      STATE_F: begin
        if (w)
          next_state = STATE_C;
        else
          next_state = STATE_D;
      end
      default: begin
        next_state = STATE_A;
      end
    endcase
  end

  assign z = current_state;
endmodule
