
module TopModule (
  input [3:0] in,
  output [2:0] out_both,
  output [3:1] out_any,
  output [3:0] out_different
);
assign out_both[0] = 1'b0; // no left neighbour for bit 0
assign out_both[1] = in[0] & in[1];
assign out_both[2] = in[1] & in[2];
assign out_both[3] = in[2];

always @(posedge clk) begin
    out_any[0] = 1'b0; // no right neighbour for bit 0
    out_any[1] = (in[0] | in[1]);
    out_any[2] = (in[1] | in[2]);
    out_any[3] = (in[2] | in[3]) || (in[0]); // wrap around for bit 3
end

always @(posedge clk) begin
    out_different[0] = 1'b0; // no left neighbour for bit 0
    out_different[1] = ~(in[0] ^ in[1]);
    out_different[2] = ~(in[1] ^ in[2]);
    out_different[3] = ~(in[2] ^ in[0]); // wrap around for bit 3
end

// VERILOG-EVAL: endmodule not found
