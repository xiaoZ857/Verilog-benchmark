
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
always @(posedge clk or posedge reset) begin
  if (reset)
    current_state <= A;
  else
    case (current_state)
      A: begin
        if (w)
          next_state <= B;
        else
          next_state <= A;
      end
      B: begin
        if (w)
          next_state <= C;
        else
          next_state <= D;
      end
      C: begin
        if (w)
          next_state <= E;
        else
          next_state <= D;
      end
      D: begin
        if (w)
          next_state <= F;
        else
          next_state <= A;
      end
      E: begin
        if (!w)
          next_state <= D;
        else
          next_state <= E;
      end
      F: begin
        next_state <= C;
      enddefault:
        $display("Invalid state transition: %b", current_state);
    endcase
  assign z = (current_state == A) ? 0 : ((current_state == B) ? 1 : ((current_state == C) ? 2 : ((current_state == D) ? 3 : ((current_state == E) ? 4 : 5))));
end

// VERILOG-EVAL: endmodule not found
