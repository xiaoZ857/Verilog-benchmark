

module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  output walk_left,
  output walk_right
);

reg [1:0] state, next_state;

localparam IDLE_LEFT = 2'b00;
localparam WALK_RIGHT = 2'b01;

always @(*) begin
    case (state)
        IDLE_LEFT: begin
            if (bump_left) 
                next_state = WALK_RIGHT;
            else 
                next_state = IDLE_LEFT;
        end

        WALK_RIGHT: begin
            if (bump_right) 
                next_state = IDLE_LEFT;
            else 
                next_state = WALK_RIGHT;
        end

        default: 
            next_state = IDLE_LEFT;
    endcase
end

always @(posedge clk or posedge areset) begin
    if (areset)
        state <= IDLE_LEFT;
    else
        state <= next_state;
end

assign walk_left = (state == IDLE_LEFT);
assign walk_right = (state == WALK_RIGHT);

endmodule
