
module TopModule (
  output out
);

  // Assign 0 to the output 'out'
  out = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
