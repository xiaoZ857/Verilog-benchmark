

module TopModule (
  output zero
);

output zero = 0;
endmodule
