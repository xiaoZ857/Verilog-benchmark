
// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.
Build a combinational circuit with two inputs, a and b. There are 7
outputs, each with a logic gate driving it:

  (1) out_and: a and b
  (2) out_or: a or b
  (3) out_xor: a xor b
  (4) out_nand: a nand b
  (5) out_nor: a nor b
  (6) out_xnor: a xnor b
  (7) out_anotb: a and-not b

module TopModule (
  input a,
  input b,
  output out_and,
  output out_or,
  output out_xor,
  output out_nand,
  output out_nor,
  output out_xnor,
  output out_anotb
);

// Module body
assign out_and = a & b;
assign out_or = a | b;
assign out_xor = a ^ b;
assign out_nand = !(a & b);
assign out_nor = !(a | b);
assign out_xnor = !(a ^ b);
assign out_anotb = a & (~b);

endmodule

// VERILOG-EVAL: errant inclusion of module definition
