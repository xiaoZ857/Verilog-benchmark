

module TopModule (
  input a,
  input b,
  input c,
  output out
);



// VERILOG-EVAL: endmodule not found
