

module TopModule (
  input [7:0] in,
  output parity
);



// VERILOG-EVAL: endmodule not found
