
module TopModule (
  input [99:0] in,
  output out_and,
  output out_or,
  output out_xor
);
  // 100-input AND gate: output is 1 only if all bits are 1
  assign out_and = &in;

  // 100-input OR gate: output is 1 if at least one bit is 1
  assign out_or = |in;

  // 100-input XOR gate: output is 1 if an odd number of bits are 1
  assign out_xor = ^in;

endmodule
