
// 4‑bit wide, 256‑to‑1 multiplexer
//  in  : 1024‑bit vector containing 256 4‑bit words (in[3:0], in[7:4], …)
//  sel : 8‑bit select (0‑255)
//  out : 4‑bit output chosen by sel
module TopModule (
    input  wire [1023:0] in,
    input  wire [7:0]    sel,
    output wire [3:0]    out
);

    // Variable part‑select: start at sel*4, take 4 bits
    assign out = in[sel*4 +: 4];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
