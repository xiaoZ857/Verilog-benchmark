

module TopModule (
  input clk,
  input reset,
  input [31:0] in,
  output reg [31:0] out
);



// VERILOG-EVAL: endmodule not found
