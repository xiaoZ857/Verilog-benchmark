
module TopModule (
  input in,
  output out
);

  // Continuous assignment for combinational logic
  assign out = in;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
