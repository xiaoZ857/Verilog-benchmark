

module TopModule (
  input wire clk,
  input wire reset,
  input wire data,
  output wire [3:0] count,
  output reg counting,
  output reg done,
  input wire ack
);

reg [3:0] delay;
reg [9:0] count;
reg counting = 0;
reg done = 0;

always @(posedge clk) begin
    if (reset) begin
        delay <= 4'b0000;
        counting <= 0;
        done <= 1;
    end else if (data == 2'b11 && data[3:2] == 2'b01) begin
        delay <= 4'b1100;
        counting <= 1;
    end else if (delay != 4'b0000) begin
        count <= {delay[3:0], count};
        if (count[9:8] == 2'b00) begin
            counting <= 1;
        end else if (count[9:8] == 2'b01) begin
            counting <= 0;
            done <= 1;
        end else if (count[9:8] == 2'b10) begin
            counting <= count[7:6];
        end else if (count[9:8] == 2'b11) begin
            counting <= count[5:4];
        end
    end
end

assign done = counting;
assign count = counting ? {delay[3:0], count[9:8]} : 10'b111111111;

always @(posedge clk or ack) begin
    if (ack && !done) begin
        delay <= 4'b0000;
        counting <= 0;
    end
end

assign counting = ~done;

// VERILOG-EVAL: endmodule not found
