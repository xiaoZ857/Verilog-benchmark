
module TopModule (
  input in1,
  input in2,
  input in3,
  output logic out
);


// VERILOG-EVAL: endmodule not found
