

module TopModule (
  input in,
  output out
);



// VERILOG-EVAL: endmodule not found
