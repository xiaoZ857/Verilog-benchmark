

module TopModule (
  input [4:1] x,
  output logic f
);



// VERILOG-EVAL: endmodule not found
