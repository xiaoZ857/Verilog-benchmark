

module TopModule (
  input clk,
  input a,
  output reg [2:0] q
);



// VERILOG-EVAL: endmodule not found
