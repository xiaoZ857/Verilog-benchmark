
`timescale 1ns / 1ps

module TopModule (
    input  wire        clk,    // Positive‑edge clock
    input  wire        reset,  // Active‑high synchronous reset
    output reg  [3:0]  q       // 4‑bit counter output
);

    // ------------------------------------------------------------------
    // Parameters
    // ------------------------------------------------------------------
    localparam MAX_COUNT = 4'd10;   // Highest value before wrap‑around

    // ------------------------------------------------------------------
    // Sequential logic – synchronous counter
    // ------------------------------------------------------------------
    always @(posedge clk) begin
        if (reset) begin
            // Reset the counter to 1
            q <= 4'd1;
        end
        else if (q == MAX_COUNT) begin
            // Wrap‑around: after 10 go back to 1
            q <= 4'd1;
        end
        else begin
            // Normal increment
            q <= q + 1'b1;
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
