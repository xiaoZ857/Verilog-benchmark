
module TopModule (
  input clk,
  input [7:0] d,
  output reg [7:0] q
);

  // Instantiate 8 D flip-flops
  reg [0:0] ff0;
  reg [0:0] ff1;
  reg [0:0] ff2;
  reg [0:0] ff3;
  reg [0:0] ff4;
  reg [0:0] ff5;
  reg [0:0] ff6;
  reg [0:0] ff7;

  always @(posedge clk) begin
    q[0] <= d[0];
    q[1] <= d[1];
    q[2] <= d[2];
    q[3] <= d[3];
    q[4] <= d[4];
    q[5] <= d[5];
    q[6] <= d[6];
    q[7] <= d[7];
  end

endmodule

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
