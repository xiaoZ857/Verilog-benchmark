
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);

reg [1:0] state;
reg [7:0] byte1, byte2, byte3;
reg done_reg;

parameter IDLE = 2'b00;
parameter BYTE1 = 2'b01;
parameter BYTE2 = 2'b10;

always @(posedge clk) begin
  if (reset) begin
    state <= IDLE;
    done_reg <= 1'b0;
    byte1 <= 8'b0;
    byte2 <= 8'b0;
    byte3 <= 8'b0;
  end else begin
    case (state)
      IDLE: begin
        done_reg <= 1'b0;
        if (in[3]) begin
          byte1 <= in;
          state <= BYTE1;
        end
      end
      
      BYTE1: begin
        byte2 <= in;
        state <= BYTE2;
      end
      
      BYTE2: begin
        byte3 <= in;
        done_reg <= 1'b1;
        state <= IDLE;
      end
      
      default: begin
        state <= IDLE;
      end
    endcase
  end
end

assign done = done_reg;
assign out_bytes = {byte1, byte2, byte3};

endmodule
