
module TopModule (
  input wire clk,
  input wire reset,
  input wire data,
  output wire [3:0] count,
  output reg counting,
  output reg done,
  input wire ack
);
reg [3:0] state;
reg [3:0] shift_reg;
reg [3:0] delay;
reg [19:0] counter;
wire [3:0] current_count;

assign count = (counting) ? 20'b1111_1111_1111_1111_0000 - counter[15:0] : 4'bxxxx;
assign current_count = counting ? 4'd10 - counter[19:16] : 4'bxxxx;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        state <= 4'd0;
        shift_reg <= 4'b0000;
        delay <= 4'b0000;
        counting <= 1'b0;
        done <= 1'b0;
        counter <= 20'd0;
    end else begin
        case (state)
            4'd0: // Detect start pattern 1101
                if (shift_reg == 4'b1101) begin
                    state <= 4'd1;
                end else begin
                    shift_reg <= {shift_reg[2:0], data};
                end
            4'd1: // Shift in duration bits
                if (counter < 20'd1000) begin
                    counter <= counter + 1;
                    if (counter == 20'd999) begin
                        delay <= {delay[2:0], data};
                        if (shift_reg == 4'b1111) begin
                            state <= 4'd2;
                            counting <= 1'b1;
                            counter <= 20'd0;
                        end
                    end
                end
            4'd2: // Counting period
                if (counter < (delay + 4'd1) * 20'd1000) begin
                    counter <= counter + 1;
                end else begin
                    state <= 4'd3;
                    counting <= 1'b0;
                    done <= 1'b1;
                end
            4'd3: // Wait for acknowledgment
                if (ack == 1'b1) begin
                    state <= 4'd0;
                    shift_reg <= 4'b0000;
                    delay <= 4'b0000;
                    done <= 1'b0;
                end
        endcase
    end
end

endmodule
