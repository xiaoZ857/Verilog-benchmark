
module TopModule (
  input [4:1] x,
  output logic f
);
always @(posedge clk) begin
    casex(x)
        3'b000 : f = 0;
        3'b001 : f = 1'b0;
        3'b110 : f = 1'b1;
        3'b111 : f = 1'b1;
        4'b0101 : f = 1'b0;
        4'b1011 : f = 1'b1;
        4'b1101 : f = 1'b1;
        4'b1110 : f = 1'b0;
        default : f = 1'bx; // x represents don't care in Karnaugh map
    endcase
end
endmodule
