
module TopModule (
  input wire clk,
  input wire reset,
  input wire data,
  output wire [3:0] count,
  output reg counting,
  output reg done,
  input wire ack
);
always @(posedge clk) begin
    if (reset) begin
        state <= IDLE;
        shift_reg <= 4'b0;
        bit_count <= 2'b0;
        delay <= 4'b0;
        timer <= 10'b0;
        counting <= 1'b0;
        done <= 1'b0;
    end else begin
        case (state)
            IDLE: begin
                shift_reg <= {shift_reg[2:0], data};
                if (shift_reg == 4'b1101) begin
                    state <= READ_DELAY;
                    bit_count <= 2'b0;
                end
                counting <= 1'b0;
                done <= 1'b0;
            end
            READ_DELAY: begin
                delay <= {delay[2:0], data};
                bit_count <= bit_count + 1;
                if (bit_count == 2'b11) begin
                    state <= COUNTING;
                    timer <= 10'd1000;
                end
                counting <= 1'b0;
                done <= 1'b0;
            end
            COUNTING: begin
                counting <= 1'b1;
                done <= 1'b0;
                if (timer > 1) begin
                    timer <= timer - 1;
                end else begin
                    timer <= 10'd1000;
                    if (delay > 0) begin
                        delay <= delay - 1;
                    end else begin
                        state <= DONE;
                        counting <= 1'b0;
                    end
                end
            end
            DONE: begin
                done <= 1'b1;
                counting <= 1'b0;
                if (ack) begin
                    state <= IDLE;
                    shift_reg <= 4'b0;
                end
            end
            default: state <= IDLE;
        endcase
    end
end

assign count = (state == COUNTING) ? delay : 4'b0;

localparam IDLE = 2'b00,
           READ_DELAY = 2'b01,
           COUNTING = 2'b10,
           DONE = 2'b11;

reg [1:0] state;
reg [3:0] shift_reg;
reg [1:0] bit_count;
reg [3:0] delay;
reg [9:0] timer;

endmodule
