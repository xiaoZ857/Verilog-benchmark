
module TopModule (
  input clk,
  input a,
  output reg [2:0] q

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
