
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output q
);
q = b OR c

// VERILOG-EVAL: endmodule not found
