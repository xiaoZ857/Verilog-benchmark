
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);
// State machine to detect PS/2 mouse protocol message boundaries
localparam IDLE = 2'b00;  // Looking for byte 1 (in[3]=1)
localparam BYTE2 = 2'b01; // Found byte 1, receiving byte 2
localparam BYTE3 = 2'b10; // Found byte 2, receiving byte 3

reg [1:0] state, next_state;

// State transition logic
always @(posedge clk) begin
  if (reset) begin
    state <= IDLE;
  end else begin
    state <= next_state;
  end
end

// Next state and output logic
always @(*) begin
  // Default values
  next_state = state;
  done = 1'b0;
  
  case (state)
    IDLE: begin
      // Wait for byte with in[3]=1 (potential start of message)
      if (in[3]) begin
        next_state = BYTE2;
      end
    end
    
    BYTE2: begin
      // We've received byte 1 in previous cycle, now receiving byte 2
      // Move to BYTE3 state for next byte
      next_state = BYTE3;
    end
    
    BYTE3: begin
      // We've received byte 2 in previous cycle, now receiving byte 3
      // Signal done since we've received all 3 bytes
      done = 1'b1;
      // Check if this byte (byte 3) could be start of next message
      if (in[3]) begin
        next_state = BYTE2;
      end else begin
        next_state = IDLE;
      end
    end
  endcase
end

// VERILOG-EVAL: endmodule not found
