
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output reg walk_left,
  output reg walk_right,
  output reg aaah,
  output reg digging
);

reg state, prev_ground;
always @(posedge clk) begin
  if (areset) begin
    state <= 0; // Reset to walking left
  end
  else begin
    case (state)
      0: begin
        if (ground) begin
          state <= 1; // Start digging if ground and dig is set
        end
        else if (bump_left || bump_right) begin
          state <= 2'b10; // Change direction if bumped
        end
      end,
      1: begin
        if (!ground && !aaah) begin // Falling
          aaah <= 1;
        end
        else if (digging) begin // Digging
          state <= 3; // Keep digging until ground is gone
        end
        else if (bump_left || bump_right) begin // Bumped while walking or falling
          // No change in direction
        end
      end,
      2: begin
        if (ground) begin
          state <= 0; // Switch to walking right
        end
        else if (!aaah && !digging) begin // Being bumped while not walking or digging
          state <= 2'b10; // Change direction
        end
      end,
      3: begin
        if (ground) begin
          state <= 0; // Stop digging and resume walking once ground is back
        end
      end
    endcase

    prev_ground <= ground;
    walk_left <= state == 0;
    walk_right <= state == 2'b10;
    digging <= state == 1 || state == 3;
    aaah <= state == 1 && !prev_ground && !digging;
  end
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
