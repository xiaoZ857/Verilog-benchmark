
module TopModule (
  input [2:0] a,
  output reg [15:0] q
);
always @* begin
    if(a[2] == 3) q <= 5a0e;
    else if(a[2] == 1 && a[1] == ee) q <= aee0;
    else if(a[2] == 2) q <= 27d4;
    else if(a[2] == 0 && a[1] == 3) q <= 1232;
    else if(a[2] == 5) q <= 64ce;
    else if(a[2] == 6 && a[1] == 5) q <= c526;
    else if(a[2] == 7) q <= 2f19;
    else q <= 0;
end

// VERILOG-EVAL: endmodule not found
