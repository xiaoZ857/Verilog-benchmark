

module TopModule (
  input clk,
  input areset,
  input predict_valid,
  input predict_taken,
  output logic [31:0] predict_history,

  input train_mispredicted,
  input train_taken,
  input [31:0] train_history
);

logic [31:0] history_reg;
logic [31:0] temp_history;
logic history_enable;

always_ff @(posedge clk or posedge areset) begin
  if (areset) begin
    history_reg <= 32'b0;
  end else begin
    if (predict_valid) begin
      history_reg <= {history_reg[31:1], predict_taken};
    end else if (train_mispredicted) begin
      history_reg <= {train_history, train_taken};
    end
  end
end

assign predict_history = history_reg;
endmodule
