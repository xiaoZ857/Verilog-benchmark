
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  output walk_left,
  output walk_right,
  output aaah
);
  reg [1:0] state, next_state;
  parameter WL = 2'b00, WR = 2'b01, FL = 2'b10, FR = 2'b11;
  
  // State register
  always @(posedge clk, posedge areset) begin
    if (areset)
      state <= WL;
    else
      state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      WL: begin
        if (~ground)
          next_state = FL;
        else if (bump_left)
          next_state = WR;
        else
          next_state = WL;
      end
      WR: begin
        if (~ground)
          next_state = FR;
        else if (bump_right)
          next_state = WL;
        else
          next_state = WR;
      end
      FL: begin
        if (ground)
          next_state = WL;
        else
          next_state = FL;
      end
      FR: begin
        if (ground)
          next_state = WR;
        else
          next_state = FR;
      end
      default: next_state = WL;
    endcase
  end
  
  // Output logic (Moore)
  assign walk_left = (state == WL);
  assign walk_right = (state == WR);
  assign aaah = state[1];
endmodule
