
module TopModule (
  input [4:1] x,
  output logic f
);

// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.
Consider the function f shown in the Karnaugh map below. d is don't-care,
which means you may choose to output whatever value is convenient.
Implement this function.

                x[1]x[2]
  x[3]x[4]   00

// VERILOG-EVAL: endmodule not found
