
module TopModule (
  input a,
  input b,
  output out_assign,
  output reg out_alwaysblock
);

  // AND gate using assign statement
  assign out_assign = a & b;

  // AND gate using combinational always block
  always @(a, b) begin
    out_alwaysblock = a & b;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
