
module TopModule (
  input a,
  input b,
  output out
);


// VERILOG-EVAL: endmodule not found
