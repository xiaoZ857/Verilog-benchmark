
module TopModule (
  input clk,
  input in,
  input reset,
  output done
);

reg [2:0] state;
reg [3:0] bit_count;
localparam IDLE = 3'd0;
localparam START = 3'd1;
localparam DATA = 3'd2;
localparam STOP = 3'd3;
localparam WAIT_STOP = 3'd4;

always @(posedge clk) begin
  if (reset) begin
    state <= IDLE;
    bit_count <= 4'd0;
    done <= 1'b0;
  end else begin
    case (state)
      IDLE: begin
        done <= 1'b0;
        if (in == 1'b0) begin  // Start bit detected
          state <= START;
          bit_count <= 4'd0;
        end
     

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
