
module TopModule (
  input c,
  input d,
  output [3:0] mux_in
);
  // Generate d' using a 2-to-1 mux
  wire not_d;
  assign not_d = d ? 1'b0 : 1'b1;  // This is actually a mux: select=d, input0=1, input1=0
  
  // mux_in[0] = c + d = c ? 1 : d
  assign mux_in[0] = c ? 1'b1 : d;
  
  // mux_in[1] = 0
  assign mux_in[1] = 1'b0;
  
  // mux_in[2] = c & d = c ? d : 0
  assign mux_in[2] = c ? d : 1'b0;
  
  // mux_in[3] = c + d' = c ? 1 : d'
  assign mux_in[3] = c ? 1'b1 : not_d;
endmodule
