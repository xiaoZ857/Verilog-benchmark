
module TopModule (
    input [3:0] in,
    output out_and,
    output out_or,
    output out_xor
);

    // Calculate the AND operation for all four inputs
    assign out_and = in[0] & in[1] & in[2] & in[3];

    // Calculate the OR operation for all four inputs
    assign out_or = in[0] | in[1] | in[2] | in[3];

    // Calculate the XOR operation for all four inputs
    // Note: XOR is associative and commutative, so we can chain them directly.
    assign out_xor = in[0] ^ in[1] ^ in[2] ^ in[3];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
