
module TopModule (
  input clk,
  input a,
  input b,
  output out_assign,
  output reg out_always_comb,
  output reg out_always_ff
);

  // XOR using assign statement
  assign out_assign = a ^ b;

  // XOR using combinational always block
  always @(*) begin
    out_always_comb = a ^ b;
  end

  // XOR using clocked always block (with flip-flop for output delay)
  always @(posedge clk) begin
    out_always_ff <= a ^ b;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
