

module TopModule (
  input clk,
  input [7:0] in,
  output reg [7:0] anyedge
);

always @(posedge clk) begin
  anyedge[0] = in[0] ^ in[0];
  anyedge[1] = in[1] ^ in[1];
  anyedge[2] = in[2] ^ in[2];
  anyedge[3] = in[3] ^ in[3];
  anyedge[4] = in[4] ^ in[4];
  anyedge[5] = in[5] ^ in[5];
  anyedge[6] = in[6] ^ in[6];
  anyedge[7] = in[7] ^ in[7];
endmodule
