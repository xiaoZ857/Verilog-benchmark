
module TopModule (
  input clk,
  input enable,
  input S,
  input A,
  input B,
  input C,
  output reg Z
);
// 8-bit shift register using D flip-flops
reg [7:0] Q;

// Initialize the shift register to avoid undefined behavior
initial begin
    Q = 8'b00000000; // Ensure this matches any required initial conditions for your tests
end

always @(posedge clk) begin
    if (enable) begin
        // Shift operation: MSB is shifted in first
        Q <= {S, Q[7:1]};
    end
end

// Multiplexer logic to select one of the outputs based on A, B, C
always @(*) begin
    case ({A, B, C})
        3'b000: Z = Q[0];
        3'b001: Z = Q[1];
        3'b010: Z = Q[2];
        3'b011: Z = Q[3];
        3'b100: Z = Q[4];
        3'b101: Z = Q[5];
        3'b110: Z = Q[6];
        3'b111: Z = Q[7];
        default: Z = 1'bx; // Consider setting this to a known value if undefined states are problematic
    endcase
end

endmodule
