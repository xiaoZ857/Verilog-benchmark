
module TopModule (
  input in,
  output out
);
  assign out = in;
endmodule

// VERILOG-EVAL: errant inclusion of module definition
