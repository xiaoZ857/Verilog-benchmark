
module TopModule (
  input ring,
  input vibrate_mode,
  output ringer,
  output motor
);
assign ringer = vibrate_mode == 1'b0 ? ring : 1'b0;
assign motor = vibrate_mode == 1'b1 ? 1 : 1'b0;
endmodule
