
module TopModule (
  input [3:0] in,
  output reg [1:0] pos
);
always @(*) begin
  casez (in)
    4'b1??? : pos = 2'd3;  // in[3] is 1
    4'b01?? : pos = 2'd2;  // in[2] is 1
    4'b001? : pos = 2'd1;  // in[1] is 1
    4'b0001 : pos = 2'd0;  // in[0] is 1
    default : pos = 2'd0;  // all bits are 0
  endcase
end
endmodule
