

module TopModule (
  input clk,
  input load,
  input [9:0] data,
  output tc
);

reg [9:0] counter;

always @(posedge clk) begin
    if (load) begin
        counter <= data;
    end else if (counter != 10'b0) begin
        counter <= counter - 1'b1;
    end
    // When counter is zero, it stays zero until a new load
end

assign tc = (counter == 10'b0);

endmodule
