
module TopModule (
  output out
);
assign out = 0;

// VERILOG-EVAL: endmodule not found
