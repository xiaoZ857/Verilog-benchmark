
module TopModule (
  input clk,
  input resetn,
  input x,
  input y,
  output f,
  output g
);

reg [2:0] current_state, next_state;
reg f, g;

parameter A = 3'b000;
parameter B = 3'b001;
parameter C = 3'b010;
parameter D = 3'b011;
parameter E = 3'b100;
parameter F = 3'b101;
parameter G = 3'b110;
parameter H = 3'b111;

always @(posedge clk) begin
  if (!resetn) begin
    current_state <= A;
  end else begin
    current_state <= next_state;
  end
end

always @(*) begin
  next_state = current_state;
  case (current_state)
    A: begin
      next_state = B;
    end
    B: begin
      next_state = C;
    end
    C: begin
      if (x == 1'b1) begin
        next_state = D;
      end else begin
        next_state = C;
      end
    end
    D: begin
      if (x == 1'b0) begin
        next_state = E;
      end else begin
        next_state = C;
      end
    end
    E: begin
      if (x == 1'b1) begin
        next_state = F;
      end else if (x == 1'b0) begin
        next_state = C;
      end else begin
        next_state = E;
      end
    end
    F: begin
      if (y == 1'b1) begin
        next_state = G;
      end else begin
        next_state = H;
      end
    end
    G: begin
      next_state = G;
    end
    H: begin
      next_state = H;
    end
    default: begin
      next_state = A;
    end
  endcase
end

always @(*) begin
  f = 1'b0;
  g = 1'b0;
  
  case (current_state)
    A: begin
      f = 1'b0;
      g = 1'b0;
    end
    B: begin
      f = 1'b1;
      g = 1'b0;
    end
    C, D, E: begin
      f = 1'b0;
      g = 1'b0;
    end
    F: begin

// VERILOG-EVAL: endmodule not found
