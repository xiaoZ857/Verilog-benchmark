
module TopModule (
  input [5:0] y,
  input w,
  output reg Y1,
  output reg Y3
);

always @(posedge w) begin
  case (y)
    2'b00 : Y1 <= 1'b0; Y3 <= 1'b0;
    2'b01 : Y1 <= 1'b1; Y3 <= 1'b0;
    2'b10 : Y1 <= y[0]; Y3 <= 1'b0;
    2'b110 : Y1 <= y[2]; Y3 <= 1'b1;
    2'b111 : Y1 <= y[4]; Y3 <= y[2];
    default : Y1 <= 1'b0; Y3 <= 1'b0;
  endcase
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
