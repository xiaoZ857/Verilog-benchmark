
module TopModule (
    input  wire clk,          // system clock
    input  wire reset,        // active‑high synchronous reset
    input  wire data

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
