
module TopModule (
  input clk,
  input shift_ena,
  input count_ena,
  input data,
  output reg [3:0] q
);
always @(posedge clk) begin
    if (shift_ena)
        q <= {data, q[2:0]};
    else if (count_ena)
        q <= q - 1;
end

endmodule
