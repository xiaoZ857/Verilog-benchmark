
module TopModule (
  input clk,
  input areset,
  input load,
  input ena,
  input [3:0] data,
  output reg [3:0] q
);
always @(posedge clk) begin
    if (areset)
        q <= 4'b0;
    else if (load)
        q <= data;
    else if (ena)
        q <= {q[2:0], 1'b0};
end
endmodule
