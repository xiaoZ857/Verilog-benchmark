
module TopModule (
  input clk,
  input reset,
  output reg [3:0] q
);

always @(posedge clk) begin
    if (reset)
        q <= 4'b0001;
    else if (q == 4'b1010)  // when count reaches 10
        q <= 4'b0001;        // wrap around to 1
    else
        q <= q + 1;          // increment counter
end
endmodule
