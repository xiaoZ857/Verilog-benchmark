
module TopModule (
  input clk,
  input [7:0] d,
  input areset,
  output reg [7:0] q
);
reg [7:0] q;

always @(posedge clk) begin
    if (areset)
        q <= {8{1'b0}}; // Reset all bits to 0
    else
        q <= d;          // Load data from d
end

endmodule
