

module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);

always @(posedge clk) begin
    if (reset) begin
        q <= 1'b1;
    end else begin
        q[4] <= q[3];
        q[3] <= q[2];
        q[2] <= q[1];
        q[1] <= q[0] ^ q[5];
        q[0] <= q[5];
    end
end

assign q[5] = 1'b0;

// VERILOG-EVAL: endmodule not found
