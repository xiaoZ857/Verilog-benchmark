
// Priority Encoder Module

module TopModule (
  input [3:0] in,  // Input is a 4-bit vector (0000 to 1111)
  output reg [1:0] pos    // Output is a 2-bit vector representing the position of the first 1 bit
);

reg [3:0] bits;   // Internal reg to store input bits

assign bits = in;

// Logic for Priority Encoder
always @(*)
begin
  if (bits[3] == 1) pos = 2'b01;  // If most significant bit is high, output is 01
  else if (bits[2] == 1 && bits[0] != 1) pos = 2'b10;  // Next bit from MSB that is not zero
  else if (bits[1] == 1 && bits[0] != 1) pos = 2'b11;  // Last non-zero bit from MSB
  else if (bits[0] == 1) pos = 2'b00;  // If all but one bit are zero, output is 00
  else pos = 2'b00;  // Output 00 for input of zeros
  
end

// Testbench Example
module TopModule TB;
  reg [3:0] in;
  reg [1:0] pos;
  
  initial begin
    in = 4'b0000;  // Start with zeros
    $dump init "Position is: pos=2'b00";
    #1000
    in = 4'b1010;
    $dump "Position is: pos=2'b10";
    #1000
    in = 4'b1101;
    $dump "Position is: pos=2'b11";
    #1000
    in = 4'b0011;
    $dump "Position is: pos=2'b01";
    #1000
    
    #5000;
    $finish;
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
