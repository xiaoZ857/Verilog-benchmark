
module TopModule (
  input clk,
  input in,
  input reset,
  output out
);


// VERILOG-EVAL: endmodule not found
