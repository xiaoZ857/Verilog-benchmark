
module TopModule (
  input clk,
  input x,
  input [2:0] y,
  output reg Y0,
  output reg z
);
reg [2:0] Y_next;
assign Y[0] = Y_next[0];

always @(posedge clk) begin
    if (x == 1'b0)
        Y_next <= y; // X=0: Next state same as present state
    else
        case(y)
            3'b000: Y_next <= 3'b001;
            3'b001: Y_next <= 3'b100;
            3'b010: Y_next <= 3'b001;
            3'b011: Y_next <= 3'b010;
            3'b100: Y_next <= 3'b100; // X=1: Next state as per table
            default: Y_next <= 3'bxxx; // Handle unexpected states
        endcase

    // Update outputs based on next state logic and condition from table
    if (Y_next == 3'b001 || Y_next == 3'b010)
        z = 1'b0;
    else if (Y_next == 3'b011 || Y_next == 3'b100)
        z = 1'b1;
end

always @(posedge clk) begin
    Y0 <= Y_next[0]; // Sequential logic for the output register
end

endmodule
