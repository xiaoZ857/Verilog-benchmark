
module TopModule (
  input [3:0] in,
  output out_and,
  output out_or,
  output out_xor
);

  // Implementing the 4-input AND gate for out_and
  assign out_and = in[0] & in[1] & in[2] & in[3];

  // Implementing the 4-input OR gate for out_or
  assign out_or = in[0] | in[1] | in[2] | in[3];

  // Implementing the 4-input XOR gate for out_xor
  // Note: A simple way to implement a 4-input XOR is by chaining two 2-input XOR gates.
  wire xor_step1, xor_step2;

  assign xor_step1 = in[0] ^ in[1];
  assign xor_step2 = in[2] ^ in[3];
  assign out_xor = xor_step1 ^ xor_step2;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
