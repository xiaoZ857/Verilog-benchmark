
module TopModule (
  input [7:0] a,
  input [7:0] b,
  output [7:0] s,
  output overflow
);
// Calculate sum using arithmetic logic units (ALUs)
logic [7:0] sum_unsigned;
assign sum_unsigned = a + b;

// Convert the sum back to its 2's complement representation
wire s_2s;
assign s_2s = ~sum_unsigned | 1; // Use bitwise OR instead of addition

// Assign the output values
assign s = s_2s[7:0];
assign overflow = (s_2s[0] == 1) && (s_2s[7] == 1);

endmodule
