
module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);

  // State encoding with 3 states
  parameter S0 = 2'b

// VERILOG-EVAL: endmodule not found
