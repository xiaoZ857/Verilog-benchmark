
assign out_xor = a ^ b; // Direct XOR operation

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
