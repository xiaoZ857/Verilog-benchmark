
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output reg out
);


// VERILOG-EVAL: endmodule not found
