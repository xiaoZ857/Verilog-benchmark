
output Y1 = (~w & y[5]) | (w & y[4]);
output Y3 = (~w & y[0]) | (w & ~y[2]);

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
