

module TopModule (
  input in,
  input [1:0] state,
  output reg [1:0] next_state,
  output out
);



// VERILOG-EVAL: endmodule not found
