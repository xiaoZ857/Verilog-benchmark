
module TopModule (
  input in,
  output out
);

  // Continuous assignment: Connect input directly to output
  assign out = in;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
