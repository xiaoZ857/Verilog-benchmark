
module TopModule (
  input c,
  input d,
  output [3:0] mux_in
);
assign mux_in[3] = a & b;
assign mux_in[2] = a | b;
assign mux_in[1] = ~a & ~b;
assign mux_in[0] = a & ~b;

endmodule
