
module TopModule (
  input in,
  input [3:0] state,
  output reg [3:0] next_state,
  output out
);

  always @(*) begin
    // State transition logic for one-hot encoding
    next_state[0] = (state[0] & ~in) | (state[2] & ~in);  // To state A
    next_state[1] = (state[0] & in) | (state[1] & in) | (state[3] & in);  // To state B
    next_state[2] = (state[1] & ~in) | (state[3] & ~in);  // To state C
    next_state[3] = state[2] & in;  // To state D
  end
  
  // Output logic (Moore machine - output depends only on current state)
  assign out = state[3];  // Output is 1 only in state D

endmodule
