
module TopModule (
  input clk,
  input a,
  input b,
  output q,
  output state
);
reg q_reg; // Register to hold the current state of q

always @(posedge clk) begin
    reg q_next; // Next state for q

    // Determine next state of q based on current inputs and state
    if (a == 1 && b == x) begin
        q_next = ~q_reg; // Toggle q when a is 1, b is don't care
    end else if (a == 0 && b == 1) begin
        q_next = 1'b1; // Set q to 1 when a is 0 and b is 1
    end else if (a == 1 && b == 1) begin
        q_next = ~q_reg; // Toggle q when both a and b are 1
    end else begin
        q_next = q_reg; // If a == 0 and b == 0, do nothing (q remains unchanged)
    end

    // Update the register holding q's value
    q_reg <= q_next;

    // Always update state to reflect current q_reg value
    state <= q_reg;
end

// Output assignment
assign q = q_reg;

endmodule
