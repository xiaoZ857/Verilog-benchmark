
module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);
assign q[0] = (q[1] ^ q[2]) & (q[3] ^ q[4]);
assign q[1] = (q[2] ^ q[3]) & (q[4] ^ q[5]);
assign q[2] = (q[3] ^ q[4]) & (q[5] ^ q[6]);
assign q[3] = (q[4] ^ q[5]) & (q[6] ^ q[7]);
assign q[4] = (q[5] ^ q[6]) & (q[7] ^ q[8]);

always @(posedge clk) begin
    if (reset)
        q <= 1'b0;
    else
        q <= {q[4], q[3], q[2], q[1], q[0]};
endmodule
