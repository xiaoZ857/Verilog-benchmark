
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out
);


// VERILOG-EVAL: endmodule not found
