
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out
);
assign out = (!a & b) | (a & !b) | (!c & d) | (c & !d);

// VERILOG-EVAL: abnormal backticks count
