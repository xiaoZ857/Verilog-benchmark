
module TopModule (
  input clk,
  input aresetn,
  input x,
  output reg z
);
// Define states using localparam
localparam S0 = 2'b00, // No bits matched
           S1 = 2'b01, // First bit '1' matched
           S2 = 2'b10; // "10" matched, waiting for '1'

reg [1:0] state, next_state;

// State register with negative edge asynchronous reset
always @(negedge clk or negedge aresetn) begin
    if (!aresetn)
        state <= S0;
    else
        state <= next_state;
end

// Next state logic (combinational)
always @(*) begin
    case (state)
        S0: next_state = x ? S1 : S0;
        S1: next_state = x ? S1 : S2;
        S2: next_state = x ? S1 : S0;
        default: next_state = S0;
    endcase
end

// Output logic (Mealy: depends on state and input)
always @(*) begin
    case (state)
        S0: z = 1'b0;
        S1: z = 1'b0;
        S2: z = x ? 1'b1 : 1'b0; // Output 1 only if current input x is '1'
        default: z = 1'b0;
    endcase
end

endmodule
