
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);
logic state;
logic next_state;

always @(posedge clk or posedge areset) begin
  if (areset) begin
    state <= 0;
  else begin
    state <= next_state;
  end
end

always @(*) begin
  case (state)
    0: begin
      if (x == 0)
        next_state = 0;
      else
        next_state = 1;
    end
    1: begin
      if (x == 0)
        next_state = 1;
      else
        next_state = 1;
    end
    default: begin
      next_state = 0;
    end
  endcase
end

assign z = state == 0 ? 0 : 1;
endmodule
