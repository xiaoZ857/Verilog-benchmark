
module TopModule (
  input clk,
  input w,
  input R,
  input E,
  input L,
  output reg Q
);


// VERILOG-EVAL: endmodule not found
