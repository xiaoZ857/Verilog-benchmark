
// Assign 0 to the output 'zero' continuously
module TopModule (
  output zero
);
  assign zero = 0;
endmodule

// VERILOG-EVAL: errant inclusion of module definition
