

module TopModule (
  input clk,
  input j,
  input k,
  output reg Q
);



// VERILOG-EVAL: endmodule not found
