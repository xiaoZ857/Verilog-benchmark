
time    a    b    q
0ns     0    0    0
5ns     0    0    0
10ns    0    0    0
15ns    0    0    0
20ns    0    0    0
25ns    0    1    0
30ns    0    1    0
35ns    1    0    0
40ns    1    0    0
45ns    1    1    1
50ns    1    1    1
55ns    0    0    0
60ns    0    0    0
65ns    0    1    0
70ns    0    1    0
75ns    1    0    0
80ns    1    0    0
85ns    1    1    1
90ns    1    1    1

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
