
module TopModule (
  input clk,
  input x,
  input [2:0] y,
  output reg Y0,
  output reg z
);
always @(posedge clk) begin
    case (y)
        3'b000: begin
            if (x) begin
                Y0 <= 1'b1;
            end else begin
                Y0 <= 1'b0;
            end
            z <= 1'b0;
        end
        3'b001: begin
            if (x) begin
                Y0 <= 1'b0;
            end else begin
                Y0 <= 1'b1;
            end
            z <= 1'b0;
        end
        3'b010: begin
            if (x) begin
                Y0 <= 1'b1;
            end else begin
                Y0 <= 1'b0;
            end
            z <= 1'b0;
        end
        3'b011: begin
            if (x) begin
                Y0 <= 1'b0;
            end else begin
                Y0 <= 1'b1;
            end
            z <= 1'b1;
        end
        3'b100: begin
            if (x) begin
                Y0 <= 1'b0;
            end else begin
                Y0 <= 1'b1;
            end
            z <= 1'b1;
        end
        default: begin
            Y0 <= 1'b0;
            z <= 1'b0;
        end
    endcase
end
endmodule
