
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output out_sop,
  output out_pos
);


// VERILOG-EVAL: endmodule not found
