
module TopModule (
  input ring,
  input vibrate_mode,
  output ringer,
  output motor
);


// VERILOG-EVAL: endmodule not found
