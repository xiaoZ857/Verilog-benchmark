
module TopModule (
  input clk,
  input shift_ena,
  input count_ena,
  input data,
  output reg [3:0] q
);

  always @(posedge clk) begin
    if (shift_ena) begin
      // Shift register: MSB first
      q[3] <= data;
      for (integer i = 3; i > 0; i--) begin
        q[i] <= q[i-1];
      end
      q[0] <= 0; // Default to 0 for the least significant bit
    end else if (count_ena) begin
      // Down counter
      q <= q - 1;
    end else begin
      // Hold the current value
      // This handles the case where neither shift_ena nor count_ena is asserted.
      // It is also important for initialization.
    end
  end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
