

module TopModule (
  input clk,
  input a,
  output reg [2:0] q
);

always @(posedge clk) begin
    if (a == 1'b1)
        q <= 3'd4;
    else if (q != 3'd0 && q != 3'd1)
        q <= q + 1'b1;
end

endmodule
