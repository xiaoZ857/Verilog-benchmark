
module TopModule(
    input clk,           // Positive clock/clk signal
    input j,              // J (reset)
    input k,              // K (set)
    output reg [1:0] Q   // Q is a 2-bit signal representing the state of the flip-flop
);

reg [1:0] Qold;

always @(posedge clk) begin
    if(k == 1 && j == 0) begin      // When K is high and J is low, set
        Q <= 1'b1;
    end else if(j == 1 && k == 0) begin // When J is high and K is low, reset
        Q <= 1'b0;
    end else if(k == 1 && j == 1) begin // When both K and J are high, toggle
        Q <= ~Qold;
    end else {                     // When K is low and J is low, retain current state
        Q <= Qold;
    }
end

always @(*) begin
    Qold = Q;         // Update the old state with the new state on each positive clock edge
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
