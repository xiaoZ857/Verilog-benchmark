
module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);
  reg [31:0] next_q;

  always @(posedge clk) begin
    if (reset) begin
      q <= 32'h1;
    end else begin
      q <= next_q;
    end
  end

  always @(*) begin
    next_q = q;
    next_q[31] = q[31] ^ q[0]; // Tap at position 32 (q[31])
    next_q[21] = q[21] ^ q[0]; // Tap at position 22 (q[21])
    next_q[1] = q[1] ^ q[0]; // Tap at position 2 (q[1])
    // No tap at position 1 (q[0])
  end

endmodule
