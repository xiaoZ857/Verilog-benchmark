
module TopModule (
  input clk,
  input slowena,
  input reset,
  output reg [3:0] q
);
always @(posedge clk) begin
  if (reset) begin
    q <= 0;
  end else if (!slowena && !reset) begin
    // do nothing
  end else if (slowena) begin
    q <= q + 1;
  end
end

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
