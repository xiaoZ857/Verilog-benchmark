

module TopModule (
  output one
);

always @(*) 
begin
    one = 1;
endmodule
