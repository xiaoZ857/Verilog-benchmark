

module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  output walk_left,
  output walk_right,
  output aaah
);

  reg state;
  reg walk_left_reg;
  reg walk_right_reg;
  reg aaah_reg;

  always @(posedge clk or posedge areset) begin
    if (areset) begin
      state <= 0; // Walk left initially
    end else begin
      case (state)
        0: begin // Walk left
          walk_left_reg <= 1;
          walk_right_reg <= 0;
          aaah_reg <= 0;
          if (bump_left) begin
            state <= 1;
          end else if (bump_right) begin
            state <= 1;
          end else if (ground == 0) begin
            state <= 2;
          end
        end
        1: begin // Walk right
          walk_left_reg <= 0;
          walk_right_reg <= 1;
          aaah_reg <= 0;
          if (bump_left) begin
            state <= 0;
          end else if (bump_right) begin
            state <= 0;
          end else if (ground == 0) begin
            state <= 2;
          end
        end
        2: begin // Falling
          walk_left_reg <= 0;
          walk_right_reg <= 0;
          aaah_reg <= 1;
          if (ground == 1) begin
            state <= (walk_left_reg == 1) ? 0 : 1;
          end
        end
        default: state <= 0;
      endcase
    end
  end

  assign walk_left = walk_left_reg;
  assign walk_right = walk_right_reg;
  assign aaah = aaah_reg;

endmodule
