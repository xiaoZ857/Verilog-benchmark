
module TopModule (
    input wire clk,
    input wire areset,
    input wire load,
    input wire ena,
    input wire [3:0] data,
    output reg [3:0] q
);

    // Asynchronous reset and synchronous operations
    always @(posedge clk or posedge areset) begin
        if (areset) begin
            // Reset the shift register to zero on asynchronous reset
            q <= 4'b0000;
        end else begin
            if (load) begin
                // Load data into the shift register when load is asserted
                q <= data;
            end else if (ena) begin
                // Shift right operation when enable is asserted
                q <= {1'b0, q[3:1]};
            end
        end
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
