

module TopModule (
  input x3,
  input x2,
  input x1,
  output f
);



// VERILOG-EVAL: endmodule not found
