
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  output walk_left,
  output walk_right,
  output aaah
);

// State encoding
localparam WALK_LEFT = 2'b00;
localparam WALK_RIGHT = 2'b01;
localparam FALL_LEFT = 2'b10;
localparam FALL_RIGHT = 2'b11;

reg [1:0] state, next_state;

// State transition logic
always @(*) begin
    case (state)
        WALK_LEFT: begin
            if (!ground) begin
                next_state = FALL_LEFT;
            end else if (bump_left) begin
                // Bumped on left (or both sides) → walk right
                next_state = WALK_RIGHT;
            end else if (bump_right) begin
                // Bumped on right only → walk left
                next_state = WALK_LEFT;
            end else begin
                next_state = WALK_LEFT;
            end
        end
        
        WALK_RIGHT: begin
            if (!ground) begin
                next_state = FALL_RIGHT;
            end else if (bump_right) begin
                // Bumped on right (or both sides) → walk left
                next_state = WALK_LEFT;
            end else if (bump_left) begin
                // Bumped on left only → walk right
                next_state = WALK_RIGHT;
            end else begin
                next_state = WALK_RIGHT;
            end
        end
        
        FALL_LEFT: begin
            if (ground) begin
                next_state = WALK_LEFT;
            end else begin
                next_state = FALL_LEFT;
            end
        end
        
        FALL_RIGHT: begin
            if (ground) begin
                next_state = WALK_RIGHT;
            end else begin
                next_state = FALL_RIGHT;
            end
        end
        
        default: begin
            next_state = WALK_LEFT;
        end
    endcase
end

// State update
always @(posedge clk or posedge areset) begin
    if (areset) begin
        state <= WALK_LEFT;
    end else begin
        state <= next_state;
    end
end

// Output logic (Moore machine)
assign walk_left = (state == WALK_LEFT);
assign walk_right = (state == WALK_RIGHT);
assign aaah = (state == FALL_LEFT) || (state == FALL_RIGHT);

endmodule
