
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  output walk_left,
  output walk_right
);
 ```verilog
always @(posedge clk or negedge areset) begin
    if (!areset)
        walk_left <= 1'b1;
    else if (bump_left)
        walk_left <= 0;
    else if (bump_right)
        walk_left <= 0;
    else
        walk_left <= walk_right;

    if (!areset)
        walk_right <= 1'b0;
    else if (bump_left)
        walk_right <= 1'b1;
    else if (bump_right)
        walk_right <= 0;
    else
        walk_right <= walk_left;
end

assign walk_left = walk_left_reg;
assign walk_right = walk_right_reg;

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
