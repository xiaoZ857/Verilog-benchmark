
module TopModule (
  input clk,
  input [7:0] d,
  input reset,
  output reg [7:0] q
);
always @(negedge clk) begin
  if (reset) begin
    // Synchronously reset to 0x34 on negative edge of clk
    q1 <= 4'b0011;  // Lower nibble should be '3'
    q2 <= 4'b0100;  // Upper nibble should be '4'
  end else begin
    // Capture data on the negative edge of clock when reset is not active
    q1 <= d[3:0];   // Update lower nibble with input data
    q2 <= d[7:4];   // Update upper nibble with input data
  end
end

always @(*) begin
  q = {q2, q1};     // Form the output byte by concatenating q2 and q1
end

endmodule
