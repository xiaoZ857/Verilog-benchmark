
module TopModule (
  output out
);
 ```verilog
always @* begin
    out = 0;
end
endmodule

// VERILOG-EVAL: abnormal backticks count
