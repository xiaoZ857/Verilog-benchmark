
module TopModule (
    input [2:0] clk, // input clock signal
    input [3:0] a,   // 4-bit input signal 'a'
    output reg [15:0] q // output signal 'q'
);

always @(posedge clk) begin
    if (a[1] == 0 && a[2] == 0) begin
        q <= 1232;
    end else if (a[1] == 3 && a[2] == 0) begin
        q <= 5a0e;
    end else if (a[1] == 4 && a[2] == 1) begin
        q <= 64ce;
    end else if (a[1] == 6 && a[2] == 1) begin
        q <= c526;
    end else if (a[1] == 0 && a[2] == 2) begin
        q <= 1232;
    end else if (a[1] == 3 && a[2] == 2) begin
        q <= 5a0e;
    end else if (a[1] == 6 && a[2] == 2) begin
        q <= 27d4;
    end else if (a[1] == 0 && a[2] == 3) begin
        q <= 2066;
    end else if (a[1] == 5 && a[2] == 1) begin
        q <= c526;
    end else if (a[1] == 4 && a[2] == 3) begin
        q <= 64ce;
    end else if (a[1] == 2 && a[2] == 0) begin
        q <= 27d4;
    end else 
    begin
        q <= aee0;
    end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
