
// Create 100-input AND gate
assign out_and = in[99:0];

// Create 100-input OR gate
assign out_or = ~in[0] | in[1] | in[2] | ... | in[99];

// Create 100-input XOR gate
assign out_xor = in[0] ^ in[1] ^ in[2] ^ ... ^ in[99];

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
