

module TopModule (
  input d,
  input ena,
  output logic q
);



// VERILOG-EVAL: endmodule not found
