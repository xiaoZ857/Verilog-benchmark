
module TopModule (
  output out
);

  always out = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
