
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
  // State definitions
  parameter [2:0] A = 3'b000,
                  B = 3'b001,
                  C = 3'b010,
                  D = 3'b011,
                  E = 3'b100,
                  F = 3'b101;
  
  reg [2:0] state, next_state;
  
  // State register with asynchronous reset
  always @(posedge clk or posedge reset) begin
    if (reset)
      state <= A;
    else
      state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      A: next_state = (w == 0) ? B : A;
      B: next_state = (w == 0) ? C : D;
      C: next_state = (w == 0) ? E : D;
      D: next_state = (w == 0) ? F : A;
      E: next_state = (w == 0) ? E : D;
      F: next_state = (w == 0) ? C : D;
      default: next_state = A;
    endcase
  end
  
  // Output logic - z=1 only in states E and F
  assign z = (state == E || state == F) ? 1'b1 : 1'b0;
