
module TopModule (
  input clk,
  input in,
  input reset,
  output done
);


// VERILOG-EVAL: endmodule not found
