
// TopModule.v
// ---------------------------------------------------------------
// Description:
//   A simple combinational module with no inputs.
//   The single output `out` is permanently driven to logic 0.
// ---------------------------------------------------------------
`timescale 1ns / 1ps

module TopModule (
    output out          // Single output, always 0
);

    // Continuous assignment: always drive `out` to 0
    assign out = 1'b0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
