
module TopModule (
  input [3:0] a,
  input [3:0] b,
  input [3:0] c,
  input [3:0] d,
  input [3:0] e,
  output reg [3:0] q
);
assign q = (a & b & ~c) | (~c & d & e) | (c & d & e) | (e & d);

endmodule
