
module TopModule (
  input clk,
  input reset,
  output shift_ena
);
module top_module(
    input clk,
    input reset,
    output shift_ena
);

// Initialize state variable to track shift register enable
reg shift_ena_prev = 0;

always @(posedge clk) begin
    if (reset)
        shift_ena <= 1;
    else 
        // If bit pattern is detected and shift_ena_prev is 0, set it high
        if (!shift_ena_prev && (clk == 1)) begin
            shift_ena <= 1;
            shift_ena_prev <= 1;
        end 
        // If the FSM is not in the reset state, toggle shift_ena on each clock cycle
        else if (shift_ena_prev) begin
            shift_ena <= ~shift_ena;
            shift_ena_prev <= !shift_ena;
        end 
        // In any other case, just flip-flop shift_ena to previous value
        else begin
            shift_ena <= shift_ena_prev;
            shift_ena_prev <= shift_ena;
        end
end

endmodule
