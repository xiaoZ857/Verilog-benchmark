
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output q
);
assign q = (a & ~b) | (~a & b & c) | (d & ~c);

// VERILOG-EVAL: endmodule not found
