
module TopModule (
  input clk,
  input [7:0] d,
  output reg [7:0] q
);
assign q = d;
endmodule
