
module TopModule (
    input  wire clk,
    input  wire reset,          // active‑high synchronous reset
    input  wire data,           // serial data input

    output reg  shift_ena,     

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
