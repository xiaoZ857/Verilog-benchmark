
module TopModule (
  input [5:0] y,
  input w,
  output Y1,
  output Y3
);
assign Y1 = (y[4] & ~w) | (y[2] & w);

always @(*) begin
    Y3 = (y[0] & ~w) | (y[3] & w);
end

endmodule
