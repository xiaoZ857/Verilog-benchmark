
module TopModule (
  output one
);

  assign one = 1;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
