
module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);

wire c_out;

full_adder fa0 (.a(x[0]), .b(y[0]), .c_in(1'b0), .s(sum[0]), .c_out(c_out));
full_adder fa1 (.a(x[1]), .b(y[1]), .c_in(c_out), .s(sum[1]), .c_out(c_out));
full_adder fa2 (.a(x[2]), .b(y[2]), .c_in(c_out), .s(sum[2]), .c_out(c_out));
full_adder fa3 (.a(x[3]), .b(y[3]), .c_in(c_out), .s(sum[3]), .c_out(c_out));

assign sum[4] = c_out;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
