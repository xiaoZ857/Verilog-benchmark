
module TopModule (
  input [3:0] a,
  input [3:0] b,
  input [3:0] c,
  input [3:0] d,
  input [3:0] e,
  output reg [3:0] q
);
always @(*) begin
    case (c)
        0: q = b;
        1: q = e;
        2: q = a;
        3: q = d;
        4: q = f;
        5: q = f;
        6: q = f;
        7: q = f;
        8: q = f;
        9: q = f;
        default: q = 4'b0;
    endcase
endmodule
