
module TopModule (
    input sel,
    input [7:0] a,
    input [7:0] b,
    output reg [7:0] out
);

always @(posedge clk) begin
    if(sel)
        out = b;
    else
        out = a;
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
