
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output q
);


// VERILOG-EVAL: endmodule not found
