
module TopModule (
  input clk,
  input d,
  input ar,
  output logic q
);

  logic q_internal;

  always_ff @(posedge clk, posedge ar) begin
    if (ar) begin
      q_internal <= 1'b0;
    end else begin
      q_internal <= d;
    end
  end

  assign q = q_internal;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
