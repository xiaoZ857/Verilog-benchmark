
module TopModule (
  input in,
  input [1:0] state,
  output reg [1:0] next_state,
  output out
);
always @(*) begin
    case (state)
        2'b00: begin // State A
            next_state = in ? 2'b01 : 2'b00; // A -> B if in=1, else A
        end
        2'b01: begin // State B
            next_state = in ? 2'b01 : 2'b10; // B -> B if in=1, else C
        end
        2'b10: begin // State C
            next_state = in ? 2'b11 : 2'b00; // C -> D if in=1, else A
        end
        2'b11: begin // State D
            next_state = in ? 2'b01 : 2'b10; // D -> B if in=1, else C
        end
    endcase
end

assign out = (state == 2'b11) ? 1'b1 : 1'b0;
endmodule
