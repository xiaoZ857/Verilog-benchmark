
module TopModule (
  input [99:0] in,
  output reg [99:0] out
);
 ```verilog
always @(posedge clk) begin
    for (int i = 0; i < 100; i++)
        out[i] <= in[99-i];
end

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
