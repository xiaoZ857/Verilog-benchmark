
// ---------------------------------------------------------------------------
//  TopModule
//  Recognizes the 8‑bit scancodes for the numeric keys 0‑9
//  and produces a 4‑bit key code together with a validity flag.
// ---------------------------------------------------------------------------

module TopModule (
    input  wire [7:0] code,   // 8‑bit keyboard scancode
    output reg  [3:0] out,    // 4‑bit key number (0‑9)
    output reg        valid   // 1‑bit flag: 1 if a key was recognized
);

    // ---------------------------------------------------------------
    //  Combinational logic: interpret the scancode
    // ---------------------------------------------------------------
    always @(*) begin
        // Default: no key matched
        out   = 4'd0;
        valid = 1'b0;

        case (code)
            8'h45: begin out = 4'd0; valid = 1'b1; end   // '0'
            8'h16: begin out = 4'd1; valid = 1'b1; end   // '1'
            8'h1e: begin out = 4'd2; valid = 1'b1; end   // '2'
            8'h26: begin out = 4'd3; valid = 1'b1; end   // '3'
            8'h25: begin out = 4'd4; valid = 1'b1; end   // '4'
            8'h2e: begin out = 4'd5; valid = 1'b1; end   // '5'
            8'h36: begin out = 4'd6; valid = 1'b1; end   // '6'
            8'h3d: begin out = 4'd7; valid = 1'b1; end   // '7'
            8'h3e: begin out = 4'd8; valid = 1'b1; end   // '8'
            8'h46: begin out = 4'd9; valid = 1'b1; end   // '9'
            default: begin out = 4'd0; valid = 1'b0; end // no match
        endcase
    end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
