
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);
assign out_byte = (in[7:0] == 8'b11110000) && (in[8] == 1'b1);
assign done = (in[7:0] == 8'b11110000) && (in[8] == 1'b1);

always @(posedge clk or reset) begin
    if (reset)
        out_byte <= 8'b00000000;
    else
        out_byte <= in[7:0];
end

assign done = done;

always @(*) begin
    if (out_byte != 8'b11110000) begin
        done <= 1'b0;
    end else begin
        done <= 1'b1;
    end
end

// VERILOG-EVAL: endmodule not found
