
module TopModule (
  output out
);
assign out = 1'b0; endmodule

// VERILOG-EVAL: endmodule not found
