
module TopModule (
  output out
);

  assign out = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
