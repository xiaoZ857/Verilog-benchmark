

module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);



// VERILOG-EVAL: endmodule not found
