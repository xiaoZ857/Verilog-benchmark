
module TopModule (
    input [2:0] a,
    input [2:0] b,
    output [2:0] out_or_bitwise,
    output out_or_logical,
    output [5:0] out_not
);

    // Compute the bitwise-OR of a and b
    assign out_or_bitwise = a | b;

    // Compute the logical-OR of a and b
    assign out_or_logical = |a | |b;  // '|' is the reduction OR operator

    // Compute the NOT (inverse) of both vectors
    assign out_not[5:3] = ~b;         // Inverse of b in upper half
    assign out_not[2:0] = ~a;         // Inverse of a in lower half

endmodule

// VERILOG-EVAL: errant inclusion of module definition
