
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);

reg [1:0] state;
reg [1:0] next_state;

always @(posedge clk or posedge areset) begin
    if (areset) begin
        state <= 2'b01;
    end else begin
        state <= next_state;
    end
end

always @(*) begin
    case (state)
        2'b01: begin
            if (x) begin
                next_state = 2'b10;
            end else begin
                next_state = 2'b01;
            end
        end
        2'b10: begin
            next_state = 2'b10;
        end
        default: begin
            next_state = 2'b01;
        end
    endcase
end

assign z = (state == 2'b01 && x) || (state == 2'b10 && ~x);

endmodule
