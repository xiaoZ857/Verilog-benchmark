
module TopModule (
  input clk,
  input reset,
  input w,
  output z
);
always @(posedge clk) begin
    if (reset)
        state <= 3'b000;
    else
        case (state)
            3'b000: state <= w ? 3'b000 : 3'b001;
            3'b001: state <= w ? 3'b011 : 3'b010;
            3'b010: state <= w ? 3'b011 : 3'b100;
            3'b011: state <= w ? 3'b000 : 3'b101;
            3'b100: state <= w ? 3'b011 : 3'b100;
            3'b101: state <= w ? 3'b011 : 3'b010;
            default: state <= 3'b000;
        endcase
end

assign z = (state == 3'b100) | (state == 3'b101);

endmodule
