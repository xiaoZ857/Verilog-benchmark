
module TopModule (
  input clk,
  input reset,
  output [3:1] ena,
  output reg [15:0] q
);
always @(posedge clk or posedge reset) begin
    if (reset) begin
        q <= 16'b0000_0000_0000_0000;
    end else begin
        {ena[3], q[3:0]} <= q[3:0] + 4'd1;
        
        if (q[3:0] == 4'd9) begin
            q[7:4] <= q[7:4] + 4'd1;
            ena[3] = 1'b1;
        end else begin
            ena[3] = 1'b0;
        end
        
        if (q[7:4] == 4'd9) begin
            {ena[2], q[11:8]} <= q[11:8] + 4'd1;
            
            if (q[11:8] == 4'd9) begin
                q[15:12] <= q[15:12] + 4'd1;
                ena[2] = 1'b1;
            end else begin
                ena[2] = 1'b0;
            end
        end else begin
            ena[2] = 1'b0;
        end
        
        if (q[11:8] == 4'd9) begin
            {ena[1], q[15:12]} <= q[15:12] + 4'd1;
            
            if (q[15:12] == 4'd9) begin
                ena[1] = 1'b1;
            end else begin
                ena[1] = 1'b0;
            end
        end else begin
            ena[1] = 1'b0;
        end
        
        if (q[15:12] == 4'd9) begin
            q <= 16'b0000_0000_0000_0000;
            
            ena[1] = 1'b1;
            ena[2] = 1'b1;
            ena[3] = 1'b1;
        end else begin
            ena[1] = 1'b0;
        end
    end
end

endmodule
