
module TopModule (
  input clk,
  input in,
  input reset,
  output done
);
always @(posedge clk or posedge reset) begin
    if (reset) begin
        state <= IDLE;
        done <= 1'b0;
        data_reg <= 8'b0;
        bit_counter <= 3'b0;
        start_bit_valid <= 1'b0; // Add a flag to track valid start bit
    end else begin
        case (state)
            IDLE: begin
                if (!in) begin
                    next_state <= START_BIT; // Potential start detected, move to verify it
                end else begin
                    next_state <= IDLE;
                end
                done <= 1'b0; // Ensure done is cleared in IDLE
            end
            
            START_BIT: begin
                if (!in) begin
                    start_bit_valid <= ~start_bit_valid; // Flip the flag to verify two consecutive low states
                    if (start_bit_valid) begin
                        data_reg <= 8'b0;
                        bit_counter <= 3'b0;
                        next_state <= RECEIVE_DATA;
                    end else begin
                        next_state <= IDLE; // Transition back only on invalid start signal
                    end
                end else begin
                    next_state <= IDLE; // If the line goes high, it's not a valid start
                end
            end
            
            RECEIVE_DATA: begin
                data_reg <= {data_reg[6:0], in}; // Shift new bit into least significant position
                
                if (bit_counter == 3'b111) begin
                    next_state <= STOP_BIT;
                end else begin
                    bit_counter <= bit_counter + 1'b1; // Increment the counter after each bit reception
                end
            end
            
            STOP_BIT: begin
                if (in) begin
                    done <= 1'b1; // Valid stop bit detected, signal completion
                    next_state <= IDLE;
                end else begin
                    next_state <= STOP_BIT; // Continue waiting for a valid high stop bit
                end
            end
            
        endcase

        state <= next_state; // Update the current state at the end of each cycle
    end
end

// VERILOG-EVAL: endmodule not found
