
module TopModule (
  input clk,
  input a,
  input b,
  output q,
  output state
);


// VERILOG-EVAL: endmodule not found
