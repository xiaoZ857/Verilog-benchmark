
module TopModule (
  input clk,
  input [7:0] d,
  input areset,
  output reg [7:0] q
);


// VERILOG-EVAL: endmodule not found
