
module TopModule (
  input [254:0] in,
  output reg [7:0] out
);
always @(*) begin
    integer i;
    out = 8'b0; // Initialize the output to zero

    for (i = 0; i < 255; i = i + 1) begin
        if (in[i]) begin
            out = out + 1;
        end
    end
end
endmodule
