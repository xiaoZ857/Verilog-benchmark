
module TopModule (
  input clk,
  input j,
  input k,
  output reg Q
);
always @(posedge clk) begin
  if (j == 1'b0 && k == 1'b0)
    Q <= Qold; // Q remains unchanged when J and K are both 0
  else if (j == 1'b0 && k == 1'b1)
    Q <= 1'b0; // Q becomes 0 when J is 0 and K is 1
  else if (j == 1'b1 && k == 1'b0)
    Q <= 1'b1; // Q becomes 1 when J is 1 and K is 0
  else // J and K are both 1
    Q <= ~Qold; // Q becomes the complement of Qold when J and K are both 1
end

always @(posedge clk or negedge reset) begin
  if (reset)
    Q <= 1'b0; // Reset condition
  else
    Qold <= Q; // Assign current Q value to Qold for the next clock cycle
end

// VERILOG-EVAL: endmodule not found
