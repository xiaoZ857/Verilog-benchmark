
module TopModule (
  output out
);
assign out = 0;
endmodule
