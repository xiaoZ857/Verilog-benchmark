
//-----------------------------------------------------------------------------
// 4‑bit wide, 256‑to‑1 multiplexer
// in   : 1024‑bit vector that holds 256 4‑bit words (packed)
// sel  : 8‑bit select – 0 → bits[3:0], 1 → bits[7:4], …, 255 → bits[1023:1020]
// out  : 4‑bit selected word
//-----------------------------------------------------------------------------
module TopModule (
    input  wire [1023:0] in,   // 256 × 4‑bit words
    input  wire [7:0]    sel,  // 8‑bit selector
    output wire [3:0]    out   // selected 4‑bit word
);

    // Variable part‑select: select 4 bits starting at sel*4
    assign out = in[sel * 4 +: 4];

endmodule

// VERILOG-EVAL: errant inclusion of module definition
