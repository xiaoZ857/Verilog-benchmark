
module TopModule (
  output zero
);

    // Always output low
    assign zero = 0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
