
module TopModule (
  input [7:0] in,
  output reg [7:0] out
);

always @(posedge clk) begin
  out <= {in[7], in[6], in[5], in[4], in[3], in[2], in[1], in[0]};
end

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
