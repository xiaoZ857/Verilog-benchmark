
module TopModule (
  input clk,
  input areset,

  input predict_valid,
  input [6:0] predict_pc,
  output reg predict_taken,
  output reg [6:0] predict_history,

  input train_valid,
  input train_taken,
  input train_mispredicted,
  input [6:0] train_history,
  input [6:0] train_pc,
  input train_new_pc // This signal is added to store the new PC after a misprediction, if any.
);

reg [127:0] PHT; // Pattern history table (128-entry table of two-bit saturating counters)
reg [6:0] branch_history; // 7-bit global branch history register

always @(posedge clk or negedge areset) begin
    if (!areset) begin
        PHT <= 7'b0; // Reset pattern history table to zero
        branch_history <= 7'b0; // Reset branch history register to zero
    end
end

always @(posedge clk) begin
    if (train_valid && train_mispredicted) begin
        PHT[train_pc] <= train_taken ? PHT[train_pc] + 1'b1 : PHT[train_pc]; // Update PHT based on the training outcome
        branch_history <= train_history; // Store the new history for mispredictions and recover the branch history register
    end
end

always @(posedge clk) begin
    if (predict_valid) begin
        predict_taken <= PHT[pc_to_index(predict_pc)][1]; // Predict taken or not based on the PHT
        predict_history <= pc_to_index(predict_pc); // Return the branch history register state used to make the prediction
    end
end

function [6:0] pc_to_index;
    input [6:0] pc;
    variable temp [7:0];
    variable index [6:0];
    begin
        temp <= pc ^ branch_history; // XOR the PC with the branch history register to get a 7-bit index
        for (index = 0; index < 128; index = index + 1) begin
            if (temp === index) return index; // If the index matches any of the entries in PHT, return that index
        end
        // If no match found, return the least significant entry (should be initialized to zero during reset)
        return 0;
    end
endfunction

// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
