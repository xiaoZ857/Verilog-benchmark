
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
  reg [1:0] state, next_state;
  
  assign out = (state == 2'b01) ? 1'b1 : 1'b0;

  always @(*) begin
      case(state)
          2'b00: next_state = (in) ? 2'b01 : 2'b10; // A -> A or B
          2'b01: next_state = (in) ? 2'b01 : 2'b10; // B -> B or B
          2'b10: next_state = (in) ? 2'b01 : 2'b00; // B -> A or B
          default: next_state = 2'b10;
      endcase
  end

  always @(posedge clk or posedge areset) begin
      if (areset)
          state <= 2'b10; // Asynchronous reset to state B
      else
          state <= next_state;
  end
endmodule
