
module TopModule (
  input a,
  input b,
  output q
);
assign q = (a == b);

// VERILOG-EVAL: endmodule not found
