
module TopModule (
  input clk,
  input j,
  input k,
  input areset,
  output out
);

parameter OFF = 1'b0;
parameter ON  = 1'b1;

reg state, next_state;

// State register with async reset
always @(posedge clk or posedge areset) begin
    if (areset)
        state <= OFF;
    else
        state <= next_state;
end

// Next state logic
always @(*) begin
    case (state)
        OFF: next_state = j ? ON : OFF;
        ON:  next_state = k ? OFF : ON;
        default: next_state = OFF;
    endcase
end

// Output logic (Moore machine)
assign out = state;

endmodule
