
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);
reg [3:0] state; // State machine with 5 states (4 bits) to handle serial input of arbitrary length
reg Sign_bit;   // Output sign bit as a separate signal instead of embedding it in z
output reg z;   // Output is a single bit, removing the redundant reg declaration

// Add timescale directive outside of module definition as required by Xilinx
`timescale 1ns / 1ps

always @(posedge clk or negedge areset) begin
    if (!areset) begin
        // Reset the state machine when reset is asserted
        state <= 0;
        Sign_bit <= 0;
        z <= 0;
    end else begin
        case (state)
            0: begin // Initial state, start accepting input from MSB
                if (x == 1'b1) begin
                    Sign_bit <= 1'b1; // Set the sign bit if the MSB is 1 (negative number)
                end
                state <= {state[3], x}; // Shift the current state to the left and append the input LSB
            end
            1: state <= {state[3], x}; // Accept more bits until the reset is asserted
            ... // Additional states to handle more bits if needed
            default: state <= 0; // Reset the state machine if an invalid state is encountered
        endcase
        z <= Sign_bit ^ (~state[0]); // Output the 2's complement of the input based on the sign bit and the MSB of the current state
    end
end

endmodule
