
// Define the timescale outside of any module
`timescale 1ns / 1ps

module TopModule (
  input clk,
  input areset,
  input train_valid,
  input train_taken,
  output logic [1:0] state
);

always @(posedge clk or posedge areset) begin
    if (areset) begin
        state <= 2'b01; // Reset to weakly not-taken state
    end else begin
        case ({train_valid, train_taken}) 
            2'b11: begin // Increment when both train_valid and train_taken are 1
                if (state < 2'b11) state <= state + 1;
            end
            2'b10: begin // Decrement when train_valid is 1 and train_taken is 0
                if (state > 2'b00) state <= state - 1;
            end
            default: state <= state; // No change otherwise
        endcase
    end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
