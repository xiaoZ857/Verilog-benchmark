
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);


// VERILOG-EVAL: endmodule not found
