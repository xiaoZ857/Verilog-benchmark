

module TopModule (
  input clk,
  input reset,
  input x,
  output reg z
);



// VERILOG-EVAL: endmodule not found
