
module TopModule (
  input in,
  input [3:0] state,
  output reg [3:0] next_state,
  output out
);

always @(*) begin
    case(state)
        4'b0001: begin // State A
            if (in) begin
                next_state = 4'b0010; // B
            end else begin
                next_state = 4'b0001; // A
            end
        end
        4'b0010: begin // State B
            if (in) begin
                next_state = 4'b0010; // B
            end else begin
                next_state = 4'b0100; // C
            end
        end
        4'b0100: begin // State C
            if (in) begin
                next_state = 4'b1000; // D
            end else begin
                next_state = 4'b0001; // A
            end
        end
        4'b1000: begin // State D
            if (in) begin
                next_state = 4'b0010; // B
            end else begin
                next_state = 4'b0100; // C
            end
        end
        default: next_state = 4'b0001; // Default to A
    endcase
end

assign out = state[3];
endmodule
