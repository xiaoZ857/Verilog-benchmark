
module TopModule (
  input clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);
logic state;
logic data_bit;
assign done = state == 4;
assign out_byte = data_bit[7:0];
always @(posedge clk) begin
  if (reset) begin
    state <= 0;
  end else begin
    case (state)
      0: begin
        if (!in) begin
          state <= 1;
        end
      end
      1: begin
        state <= 2;
      end
      2: begin
        data_bit[0] <= in;
        state <= 3;
      end
      3: begin
        data_bit[1] <= in;
        state <= 3;
      end
      4: begin
        data_bit[2] <= in;
        state <= 3;
      end
      5: begin
        data_bit[3] <= in;
        state <= 3;
      end
      6: begin
        data_bit[4] <= in;
        state <= 3;
      end
      7: begin
        data_bit[5] <= in;
        state <= 3;
      end
      8: begin
        data_bit[6] <= in;
        state <= 3;
      end
      9: begin
        data_bit[7] <= in;
        state <= 3;
      end
      default: state <= 0;
    endcase
  end
endmodule
