
module TopModule (
  input in,
  input [1:0] state,
  output reg [1:0] next_state,
  output out
);

always @(*) begin
  case (state)
    2'b00: begin // State A
      next_state = in ? 2'b01 : 2'b00; // in=1 -> B, in=0 -> A
    end
    2'b01: begin // State B
      next_state = in ? 2'b01 : 2'b10; // in=1 -> B, in=0 -> C
    end
    2'b10: begin // State C
      next_state = in ? 2'b11 : 2'b00; // in=1 -> D, in=0 -> A
    end
    2'b11: begin // State D
      next_state = in ? 2'b01 : 2'b10; // in=1 -> B, in=0 -> C
    end
    default: next_state = 2'b00; // Default to state A
  endcase
end

// Output logic for Moore machine (output depends only on current state)
assign out = (state == 2'b11); // Only state D has output 1

endmodule
