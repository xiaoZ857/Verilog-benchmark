
module TopModule (
  input [99:0] in,
  output out_and,
  output out_or,
  output out_xor
);
assign out_and = in[99];
assign out_or = ~(~in[99] | in[98:0]);
assign out_xor = ~((in[99] & ~in[98]) | (in[98:1] & in[0]));

// VERILOG-EVAL: endmodule not found
