
module TopModule (
  input [3:0] in,
  output [2:0] out_both,
  output [3:1] out_any,
  output [3:0] out_different
);
assign out_both[2] = in[2] & in[3];
assign out_both[1] = in[1] & in[2];
assign out_both[0] = in[0] & in[1];

assign out_any[3] = in[3] | in[2];
assign out_any[2] = in[2] | in[1];
assign out_any[1] = in[1] | in[0];
assign out_any[0] = 1'b1; // Since in[0] has no neighbour to the right

always @(*) begin
    out_different[3] = in[3] ^ in[0]; // Wrapping around: in[3]'s left is in[0]
    out_different[2] = in[2] ^ in[3];
    out_different[1] = in[1] ^ in[2];
    out_different[0] = in[0] ^ in[1];
end

endmodule
