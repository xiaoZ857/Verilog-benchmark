
module TopModule (
  input [3:1] y,
  input w,
  output reg Y2
);
always @(y w) begin
  case (y[3:1])
    4'b0000: Y2 = 1'b0;
    4'b0001: Y2 = 1'b1;
    4'b0010: Y2 = 1'b1;
    4'b0011: Y2 = 1'b1;
    4'b0100: Y2 = 1'b1;
    4'b0101: Y2 = 1'b1;
    4'b0110: Y2 = 1'b1;
    4'b0111: Y2 = 1'b1;
    4'b1000: Y2 = 1'b1;
    4'b1001: Y2 = 1'b1;
    4'b1010: Y2 = 1'b1;
    4'b1011: Y2 = 1'b1;
    4'b1100: Y2 = 1'b1;
    4'b1101: Y2 = 1'b1;
    4'b1110: Y2 = 1'b1;
    4'b1111: Y2 = 1'b1;
  endcase
endmodule
