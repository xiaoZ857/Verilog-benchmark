

module TopModule (
  input in,
  output out
);

assign out = ~in;

// VERILOG-EVAL: endmodule not found
