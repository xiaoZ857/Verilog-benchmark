
module TopModule (
  input [7:0] in,
  output [7:0] out
);
always @(posedge clk) begin
    assign temp = {in[0], in[1], in[2], in[3], in[4], in[5], in[6], in[7]}; // Store input in a temporary wire for reversing
    out = temp[7:0];                                         // Assign the reversed bit order to output
end
endmodule
