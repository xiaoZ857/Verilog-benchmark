
module TopModule (
  input a,
  input b,
  input c,
  output out
);
out = a | b;

// VERILOG-EVAL: endmodule not found
