
module TopModule (
  input clk,
  input a,
  output reg [2:0] q
);
// Initialize the internal state variable 'q'
reg [2:0] q;

// Always block to update the output signal 'q'
always @(posedge clk) begin
    if (a == 1) begin
        // If input signal 'a' is high, set the output signal 'q' to 4
        q <= 4;
    else if (a == 0) begin
        // If input signal 'a' is low, update the output signal 'q'
        case(q)
            4: q = 5;   // If current value of 'q' is 4, set it to 5
            5: q = 6;   // If current value of 'q' is 5, set it to 6
            6: q = 0;   // If current value of 'q' is 6, reset it to 0
            default: q = 1; // Otherwise, set 'q' to 1
        endcase
    end
end

// Initialize the output signal 'q'
initial begin
    q <= 1;
end

endmodule
