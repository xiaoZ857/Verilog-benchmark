
module TopModule (
  input clk,
  input in,
  input areset,
  output out
);
reg A, B;

always @(posedge clk or negedge areset) begin
  if (areset) begin
    A <= 0;
    B <= 1;
  end else if (A == B) begin
    A <= in;
  end else begin
    B <= A ^ in; // XOR operation to determine next state of B
  end
end

assign out = B;

endmodule
