
module TopModule (
  input in1,
  input in2,
  input in3,
  output logic out
);
To implement the described circuit, we'll create a module that uses an

// VERILOG-EVAL: endmodule not found
