
module TopModule (
  input [99:0] in,
  output reg [99:0] out
);
always @(posedge clk) begin
  for (int i = 0; i < 100; i++) begin
    out[i] <= in[i]; // Assign the reversed bit order to the output vector
  end
end

// If you want to use blocking assignment, uncomment the following line:
// assign out[i] = in[i];

// Add clock enable if needed (assuming clk_en is an input)
// always @(posedge clk and clk_en) begin
//   for (int i = 0; i < 100; i++) begin
//     out[i] <= in[i]; // Assign the reversed bit order to the output vector
//   end
// end
endmodule
