

module TopModule (
  input clock,
  input a,
  output reg p,
  output reg q
);



// VERILOG-EVAL: endmodule not found
