
module TopModule (
  input clk,
  input enable,
  input S,
  input A,
  input B,
  input C,
  output reg Z
);
  // 8‑bit shift register (Q[0] is MSB, Q[7] is LSB)
  reg [7:0] q;

  // Shift logic: synchronous enable
  always @(posedge clk) begin
    if (enable)
      q <= {S, q[6:0]};   // Shift left, new bit S into Q[0]
  end

  // Random‑access read (3‑to‑8 mux) – combinational
  always @(*) begin
    case ({A, B, C})
      3'b000: Z = q[0];
      3'b001: Z = q[1];
      3'b010: Z = q[2];
      3'b011: Z = q[3];
      3'b100: Z = q[4];
      3'b101: Z = q[5];
      3'b110: Z = q[6];
      3'b111: Z = q[7];
      default: Z = 1'b0;   // safety default
    endcase
  end

endmodule
