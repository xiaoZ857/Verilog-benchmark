
module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);
// Initialize the state of the shift register to all ones
reg [SHIFT_REG_BITS-1:0] initialState = { SHIFT_REG_BITS-1: 1 };

// Initialize the current state of the shift register
reg [SHIFT_REG_BITS-1:0] currentState;

// Assign the initial state to the current state
always @(posedge clk or reset)
    if (reset) 
        currentState <= initialState;
    else {
        // Calculate the next state by XORing the bits at the taps with the LSB output bit
        reg [SHIFT_REG_BITS-1:0] nextState = currentState;
        for (int i = 0; i < SHIFT_REG_BITS; i++) {
            if (TAPS[i] == 0) 
                nextState[i] = currentState[i];
            else 
                nextState[i] = ~currentState[TAPS[i]];
        }

        // Update the current state to the next state
        currentState <= nextState;
    }

// Assign the output q as the LSB of the current state
assign q = currentState[0];

// Define the number of bits in the shift register
parameter SHIFT_REG_BITS = 32;

// Define the taps for the Galois LFSR
parameter TAPS = {22, 2, 1};

endmodule
