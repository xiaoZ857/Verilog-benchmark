
module TopModule (
  input clk,
  input areset,
  input bump_left,
  input bump_right,
  input ground,
  input dig,
  output walk_left,
  output walk_right,
  output aaah,
  output digging
);

// State encoding for the Lemmings FSM
parameter WALK_LEFT = 3'b000;
parameter WALK_RIGHT = 3'b001;
parameter FALL_LEFT = 3'b010;
parameter FALL_RIGHT = 3'b011;
parameter DIG_LEFT = 3'b100;
parameter DIG_RIGHT = 3'b101;
parameter SPLATTER = 3'b110;

reg [2:0] state, next_state;
reg [4:0] fall_counter; // Counter for fall duration (up to 31 cycles)

// State transition logic
always @(*) begin
  next_state = state;
  
  case (state)
    WALK_LEFT: begin
      if (!ground) begin
        next_state = FALL_LEFT;
      end else if (dig) begin
        next_state = DIG_LEFT;
      end else if (bump_left || bump_right) begin
        next_state = WALK_RIGHT;
      end
    end
    
    WALK_RIGHT: begin
      if (!ground) begin
        next_state = FALL_RIGHT;
      end else if (dig) begin
        next_state = DIG_RIGHT;
      end else if (bump_left || bump_right) begin
        next_state = WALK_LEFT;
      end
    end
    
    FALL_LEFT: begin
      if (ground) begin
        if (fall_counter > 20) begin
          next_state = SPLATTER;
        end else begin
          next_state = WALK_LEFT;
        end
      end
    end
    
    FALL_RIGHT: begin
      if (ground) begin
        if (fall_counter > 20) begin
          next_state = SPLATTER;
        end else begin
          next_state = WALK_RIGHT;
        end
      end
    end
    
    DIG_LEFT: begin
      if (!ground) begin
        next_state = FALL_LEFT;
      end
    end
    
    DIG_RIGHT: begin
      if (!ground) begin
        next_state = FALL_RIGHT;
      end
    end
    
    SPLATTER: begin
      next_state = SPLATTER; // Stay in splatter state forever
    end
  endcase

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: endmodule not found
