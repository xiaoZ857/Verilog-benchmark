
A   – reset / waiting for s
B0  – first cycle of the 3‑cycle window
B1  – second cycle
B2  – third cycle (output decision made here)

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
