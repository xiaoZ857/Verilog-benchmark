
module TopModule (
  output zero
);
assign zero = 0;
endmodule
