
//  TopModule implements a 4‑state Moore FSM
//  with one input (in), one output (out) and a synchronous active‑high reset.
//  The state transition table is:
//
//  State | Next state (in=0) | Next state (in=1) | Output
//  -----------------------------------------------------
//  A     | A                 | B                 | 0
//  B     | C                 | B                 | 0
//  C     | A                 | D                 | 0
//  D     | C                 | B                 | 1
//
//  Reset (active high) forces the FSM back to state A.
//
//  The output is a Moore output – it depends only on the current state.

module TopModule (
    input  wire clk,    // clock
    input  wire in,     // input that drives state transitions
    input  wire reset,  // synchronous active‑high reset
    output wire out     // Moore output
);

    // ------------------------------------------------------------
    // State encoding (2‑bit)
    // ------------------------------------------------------------
    localparam [1:0] STATE_A = 2'b00,
                     STATE_B = 2'b01,
                     STATE_C = 2'b10,
                     STATE_D = 2'b11;

    // Current state register
    reg [1:0] state, next_state;

    // ------------------------------------------------------------
    // Sequential logic – state register (synchronous reset)
    // ------------------------------------------------------------
    always @(posedge clk) begin
        if (reset) begin
            state <= STATE_A;          // reset to state A
        end else begin
            state <= next_state;       // normal state transition
        end
    end

    // ------------------------------------------------------------
    // Combinational logic – next state logic
    // ------------------------------------------------------------
    always @(*) begin
        case (state)
            STATE_A: begin
                if (in == 1'b0) next_state = STATE_A;
                else            next_state = STATE_B;
            end
            STATE_B: begin
                if (in == 1'b0) next_state = STATE_C;
                else            next_state = STATE_B;
            end
            STATE_C: begin
                if (in == 1'b0) next_state = STATE_A;
                else            next_state = STATE_D;
            end
            STATE_D: begin
                if (in == 1'b0) next_state = STATE_C;
                else            next_state = STATE_B;
            end
            default: next_state = STATE_A; // safety net
        endcase
    end

    // ------------------------------------------------------------
    // Output logic – Moore output (combinational)
    // ------------------------------------------------------------
    assign out = (state == STATE_D) ? 1'b1 : 1'b0;

endmodule

// VERILOG-EVAL: errant inclusion of module definition
