
module TopModule (
    input clk,
    input slowena,
    input reset,
    output

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
