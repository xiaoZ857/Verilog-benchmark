
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);
always @(posedge clk or posedge areset) begin
    if (areset) begin
        state <= 2'b01; // State A is active
    end else begin
        case (state)
            2'b01: // State A
                if (x) begin
                    state <= 2'b10; // Transition to state B
                end
                // If x=0, stay in state A (no change needed)
            2'b10: // State B
                // No conditional transitions; always stay in B
                // (since both inputs keep it in B)
                state <= 2'b10;
            default: // Should not happen, but reset to A if it does
                state <= 2'b01;
        endcase
    end
end

// Mealy output logic: z depends on current state and input x
assign z = (state == 2'b01 && x) || (state == 2'b10 && ~x);

endmodule
