
module TopModule(
    input clk,          // Positive edge triggered clock signal
    input a,             // Input signal
    output reg q         // Output register to store state
);

reg [1:0] state;      // Internal state of 2-bit counter

always @(posedge clk) begin
    if (state == 2'b00) begin
        state = a;
        q = ~a;
    elseif (state == 2'b01 && a==0) begin
        state = 2'b10;
        q = 1'b1;
    elseif (state == 2'b01 && a==1) begin
        state = 2'b00;
        q = 1'b0;
    elseif (state == 2'b10 && a==0) begin
        state = 2'b11;
        q = 1'b1;
    elseif (state == 2'b10 && a==1) begin
        state = 2'b00;
        q = 1'b0;
    elseif (state == 2'b11) begin
        state = 2'b01;
        q = 1'b1;
    end
end

endmodule

// VERILOG-EVAL: errant inclusion of module definition
