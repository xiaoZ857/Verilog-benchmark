
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);


// VERILOG-EVAL: endmodule not found
