
module TopModule (
  output out
);
  // Assign 0 to the output continuously
  assign out = 0;
endmodule

// VERILOG-EVAL: errant inclusion of module definition
