
module TopModule (
  input clk,
  input a,
  output reg q
);
  always @(posedge clk) begin
    if (a == 0) begin
      q <= 1;
    end else begin
      q <= ~q;
    end
  end

// VERILOG-EVAL: endmodule not found
