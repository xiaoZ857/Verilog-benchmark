
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);

  reg [1:0] state, next_state;
  
  // State encoding
  localparam IDLE = 2'b00;
  localparam BYTE2 = 2'b01;
  localparam BYTE3 = 2'b10;
  
  // State register
  always @(posedge clk) begin
    if (reset)
      state <= IDLE;
    else
      state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (state)
      IDLE: begin
        if (in[3])
          next_state = BYTE2;
        else
          next_state = IDLE;
      end
      
      BYTE2: begin
        next_state = BYTE3;
      end
      
      BYTE3: begin
        if (in[3])
          next_state = BYTE2;
        else
          next_state = IDLE;
      end
      
      default: next_state = IDLE;
    endcase
  end
  
  // Output logic
  assign done = (state == BYTE3);

endmodule
