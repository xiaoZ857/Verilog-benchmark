
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output [23:0] out_bytes,
  output done
);
// Finite State Machine for message boundary detection
module fsm (
  input clk,
  input reset,
  input [7:0] in,
  output [7:3][23:16] in_bound,
  output reg done,
  output [23:0] out_bytes
);

reg [3:0][23:16] state;
reg [2:0][23:16] temp_out;
reg [7:0] last_byte;

// State machine states
const int STATE_IDLE = 0;
const int STATE_BYTE_1 = 1;
const int STATE_BYTE_2 = 2;
const int STATE BYTE_3 = 3;
const int STATE-done = 4;

// States and next state values for FSM
reg [3:0] state_next;

assign state_next[STATE_IDLE]    = STATE_BYTE_1;
assign state_next[STATE_BYTE_1]   = STATE_BYTE_2;
assign state_next[STATE_BYTE_2]   = STATE_BYTE_3;
assign state_next[STATE_BYTE_3]   = STATE-done;
assign state_next[STATE_done]     = STATE_idle;

// FSM state assignment
always @(*) begin
  case(state)
    STATE_IDLE : 
      if (in[3] == 1) begin
        state = STATE_BYTE_1;
      end else begin
        state = STATE_IDLE;
      end

    STATE_BYTE_1 : 
      if (in[2] == 1) begin
        state = STATE_BYTE_2;
      end else begin
        state = STATE_IDLE;
      end

    STATE_BYTE_2 :
      if (in[1] == 1) begin
        state = STATE_BYTE_3;
      end else begin
        state = STATE_IDLE;
      end

    STATE_BYTE_3 : 
      if (in[0] == 1) begin
        state = STATE-done;
        temp_out = {in[2:0], in[1:0]};
        last_byte = in[0];
      end else begin
        state = STATE_IDLE;
        temp_out = {in[2:0], in[1:0]};
        last_byte = in[0];
      end

    STATE_done :
      if (reset) begin
        state = STATE_IDLE;
      end else begin
        state = STATE_idle;
        done = 1;
      end
  endcase
end

// FSM output signals assignment
assign in_bound[3:0] = {last_byte[2], last_byte[1], last_byte[0], temp_out[3][2]};
assign out_bytes = temp_out;

assign done = (state == STATE-done);

endmodule

// Finite state machine for message output formatting
module datapath (
  input clk,
  input reset,
  input [7:0] in_bound,
  output reg [23:0] out_bytes,
  output reg [1:0] done
);

reg [2:0][23:16] temp_out;

always @(*) begin
  if (in_bound[3:0] == {1,0,0}) begin
    // Invalid byte order
    temp_out = {1, 0, 0};
  end else begin
    temp_out = in_bound;
  end

  out_bytes = temp_out;

  done = (in_bound[3:0] == {1,0,0});

endmodule

// Main module assignment
assign in_bound[3:0] = fsm.in_bound[3:0];
assign fsm.done = fsm.done;

module TopModule (
  input clk,
  input reset,
  input [7:0] in,
  output [23:0] out_bytes,
  output done
);

TopModule top_module (
  .clk(clk),
  .reset(reset),
  .in(in),
  .out_bytes(out_bytes),
  .done(done)
);

// VERILOG-EVAL: errant inclusion of module definition
