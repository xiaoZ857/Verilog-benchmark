
module TopModule (
  input clk,
  input a,
  output reg q
);


// VERILOG-EVAL: endmodule not found
