
module TopModule (
  input clk,
  input reset,
  output reg [4:0] q
);
module top_module(
    input  clk,         // Clock signal
    input  reset_n    , // Active-low synchronous reset (Active-high for normal operation)
    output reg [4:0] q   // Output register (maximal-length state)
);

reg [1:0][4:0] shiftreg; // Internal shiftregister

// Initial values of the shiftregister
reg [1:2][4:0] tap[5:3]; // Tap positions with their initial outputs
tap[5]  = {{1,1,0,0}, {0,1,1,0}}; // Tap 5 produces output {q0,q1} 
tap[3]  = {{0,0,1,1},   {0,0,0,1}}; // Tap 3 produces output q2

// Verilog LFSR equation
reg [1:0][4:0] next_state;
always @(posedge clk or posedge reset_n) begin
    if (reset_n == 1)
        shiftreg = (tap[5][0] ^ tap[3][1]);
    else
        // XOR each output with the corresponding input bit, except for q[4]
        shiftreg[0:2] = {tap[5][0],tap[3][0],tap[5][1]};
        shiftreg[3:4] = {shiftreg[3], shiftreg[4]};
    // Update next_state
    reg [1:0][4:0] temp = (shiftreg[2:0]);
    for(int i=5;i>=3;--i) begin
        if(i != 5)
            temp[4+i-1]=temp[4+~(tap[i][0]&1)];
        else
            temp[0]=temp[0]^tap[i-1][0];
    end
    next_state = temp;
end

// Update q output
always @*(posedge clk) begin
    $regdrop q = next_state[3:4];
end

endmodule // top_module
