
module TopModule (
  input clk,
  input x,
  input [2:0] y,
  output reg Y0,
  output reg z
);

always @(posedge clk) begin
  // Implement Y[0] based on current state and input
  case (y)
    3'b000: Y0 <= x;        // Y[0]=0 when x=0, Y[0]=1 when x=1
    3'b001: Y0 <= ~x;       // Y[0]=1 when x=0, Y[0]=0 when x=1
    3'b010: Y0 <= x;        // Y[0]=0 when x=0, Y[0]=1 when x=1
    3'b011: Y0 <= ~x;       // Y[0]=1 when x=0, Y[0]=0 when x=1
    3'b100: Y0 <= ~x;       // Y[0]=1 when x=0, Y[0]=0 when x=1
    default: Y0 <= 1'b0;    // Default case for undefined states
  endcase
  
  // Implement output z based on current state
  case (y)
    3'b000: z <= 1'b0;
    3'b001: z <= 1'b0;
    3'b010: z <= 1'b0;
    3'b011: z <= 1'b1;
    3'b100: z <= 1'b1;
    default: z <= 1'b0;     // Default case for undefined states
  endcase
end

endmodule
