
module TopModule (
  input clk,
  input reset,
  output reg [31:0] q
);
always @(posedge clk or posedge reset) begin
    if (reset)
        q <= 32'h1;
    else begin
        q[31] <= ^{q[31], q[22], q[2], q[1]};
        q[30:1] <= q[29:0];
        q[0] <= q[31];
    end
end
endmodule
