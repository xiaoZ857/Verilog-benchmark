
module TopModule (
  input [3:0] in,
  output [2:0] out_both,
  output [3:1] out_any,
  output [3:0] out_different
);
always @(posedge clk) begin
  // Initialize outputs to 0
  out_both <= 3'b000;
  out_any <= 4'b0001;
  out_different <= 4'b1110;

  // Calculate out_both
  out_both[0] <= in[0];
  for (int i = 1; i < 4; i++)
    out_both[i] <= (in[i] & in[i-1]);

  // Calculate out_any
  for (int i = 1; i < 4; i++)
    out_any[i] <= (in[i] | in[(i+1)%4]);

  // Calculate out_different
  for (int i = 1; i < 4; i++)
    out_different[i] <= (in[i] ^ in[(i-1+4)%4]);
end

// Treat the vector as wrapping around, so in[3]'s neighbour to the left is in[0].

endmodule
