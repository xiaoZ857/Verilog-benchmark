
module TopModule (
  input a,
  input b,
  input c,
  input d,
  output reg out
);
  always @(a, b, c, d) begin
    out = c | d;
  end

endmodule
