
module TopModule (
  input [3:0] x,
  input [3:0] y,
  output [4:0] sum
);
wire carry0, carry1, carry2, carry3, carry4;

assign carry0 = 1'b0;
assign sum[0] = x[0] ^ y[0] ^ carry0;
assign carry1 = (x[0] & y[0]) | (carry0 & (x[0] ^ y[0]));
assign sum[1] = x[1] ^ y[1] ^ carry1;
assign carry2 = (x[1] & y[1]) | (carry1 & (x[1] ^ y[1]));
assign sum[2] = x[2] ^ y[2] ^ carry2;
assign carry3 = (x[2] & y[2]) | (carry2 & (x[2] ^ y[2]));
assign sum[3] = x[3] ^ y[3] ^ carry3;
assign carry4 = (x[3] & y[3]) | (carry3 & (x[3] ^ y[3]));
assign sum[4] = carry4;

endmodule
