

module TopModule (
  input clk,
  input reset,
  output shift_ena
);



// VERILOG-EVAL: endmodule not found
