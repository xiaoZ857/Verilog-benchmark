

module TopModule (
  input [7:0] in,
  output reg [2:0] pos
);



// VERILOG-EVAL: endmodule not found
