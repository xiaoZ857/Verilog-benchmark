
// Implement the Verilog module based on the following description. Assume that signals are positive clock/clk triggered unless otherwise stated.
Create a half adder. A half adder adds two bits (with no carry-in) and
produces a sum and carry-out.

module TopModule (
  input a,
  input b,
  output sum,
  output cout
);

  assign sum = a ^ b;  // XOR gate for sum
  assign cout = a & b; // AND gate for carry-out

endmodule

// VERILOG-EVAL: errant inclusion of module definition
