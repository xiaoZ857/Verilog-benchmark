
module TopModule (
  input clk,
  input areset,
  input x,
  output z
);

  parameter S0 = 2'b00;
  parameter S1 = 2'b01;
  parameter S2 = 2'b10;
  parameter S3 = 2'b11;
  
  reg [1:0] current_state, next_state;
  
  // State register
  always @(posedge clk or posedge areset) begin
    if (areset)
      current_state <= S0;
    else
      current_state <= next_state;
  end
  
  // Next state logic
  always @(*) begin
    case (current_state)
      S0: begin
        if (x == 0)
          next_state = S0;
        else
          next_state = S2;
      end
      S1: begin
        if (x == 0)
          next_state = S0;
        else
          next_state = S2;
      end
      S2: begin
        if (x == 0)
          next_state = S3;
        else
          next_state = S2;
      end
      S3: begin
        if (x == 0)
          next_state = S3;
        else
          next_state = S2;
      end
      default: next_state = S0;
    endcase
  end
  
  // Output logic (Moore machine - output depends only on current state)
  assign z = current_state[1];

endmodule
