
module TopModule (
  input [4:1] x,
  output logic f
);
assign f = ~x[1] & x[2];

// VERILOG-EVAL: endmodule not found
