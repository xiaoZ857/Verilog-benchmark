
module TopModule (
    input  wire clk,     // active‑high clock
    input  wire areset,  //

// VERILOG-EVAL: abnormal backticks count
// VERILOG-EVAL: errant inclusion of module definition
// VERILOG-EVAL: endmodule not found
