
module TopModule (
  input clk,
  input [7:0] in,
  input reset,
  output done
);
  always @(posedge clk) begin
    if (reset) begin
      state <= WAIT_BYTE1;
    end else begin
      state <= next_state;
    end
  end

  always @(*) begin
    case (state)
      WAIT_BYTE1: begin
        if (in[3] == 1'b1) begin
          next_state = WAIT_BYTE2;
        end else begin
          next_state = WAIT_BYTE1;
        end
      end
      WAIT_BYTE2: begin
        next_state = WAIT_BYTE3;
      end
      WAIT_BYTE3: begin
        if (in[3] == 1'b1) begin
          next_state = WAIT_BYTE2;
        end else begin
          next_state = WAIT_BYTE1;
        end
      end
      default: next_state = WAIT_BYTE1;
    endcase
  end

  assign done = (state == WAIT_BYTE3);
endmodule
