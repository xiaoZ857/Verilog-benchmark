

module TopModule (
  input clk,
  input reset,
  input data,
  output start_shifting
);

  reg [3:0] state;
  reg start_shifting_reg;

  always @(posedge clk) begin
    if (reset) begin
      state <= 0;
      start_shifting_reg <= 0;
    end else begin
      case (state)
        0: begin
          if (data == 1) begin
            state <= 1;
          end else begin
            state <= 0;
          end
        end
        1: begin
          if (data == 1) begin
            state <= 2;
          end else begin
            state <= 0;
          end
        end
        2: begin
          if (data == 0) begin
            state <= 3;
          end else begin
            state <= 0;
          end
        end
        3: begin
          if (data == 1) begin
            state <= 4;
          end else begin
            state <= 0;
          end
        end
        4: begin
          start_shifting_reg <= 1;
          state <= 4;
        end
        default: begin
          state <= 0;
        end
      endcase
    end
  end

  assign start_shifting = start_shifting_reg;
endmodule
