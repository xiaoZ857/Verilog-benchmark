
module TopModule (
  input a,
  input b,
  output out
);

// AND operation
assign out = a & b; // a AND b

endmodule

// VERILOG-EVAL: errant inclusion of module definition
